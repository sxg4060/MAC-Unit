
-- 
-- Definition of  BIST
-- 
--      Fri Dec  6 15:00:32 2019
--      
--      LeonardoSpectrum Level 3, 2008b.3
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity BIST is
   port (
      B : IN std_logic_vector (15 DOWNTO 0) ;
      C : IN std_logic_vector (15 DOWNTO 0) ;
      Cin : IN std_logic ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      test_mode : IN std_logic ;
      signature : OUT std_logic_vector (31 DOWNTO 0) ;
      mac_output : OUT std_logic_vector (31 DOWNTO 0)) ;
end BIST ;

architecture behavioral of BIST is
   signal mac_unit_tempP_31, nx1885, lfsr_C_15, test_input_lfsr_signal_15, 
      nx10, test_input_lfsr_signal_14, test_input_lfsr_signal_13, 
      test_input_lfsr_signal_12, test_input_lfsr_signal_11, 
      test_input_lfsr_signal_10, test_input_lfsr_signal_9, 
      test_input_lfsr_signal_8, test_input_lfsr_signal_7, 
      test_input_lfsr_signal_6, test_input_lfsr_signal_5, 
      test_input_lfsr_signal_4, test_input_lfsr_signal_3, 
      test_input_lfsr_signal_2, test_input_lfsr_signal_1, 
      test_input_lfsr_signal_0, nx14, nx90, nx98, lfsr_C_14, nx114, nx122, 
      lfsr_C_13, nx146, lfsr_C_12, nx170, lfsr_C_11, nx194, lfsr_C_10, nx218, 
      lfsr_C_9, nx242, lfsr_C_8, nx266, lfsr_C_7, nx290, lfsr_C_6, nx314, 
      lfsr_C_5, nx338, lfsr_C_4, nx362, lfsr_C_3, nx386, lfsr_C_2, nx410, 
      lfsr_C_1, nx434, lfsr_B_15, nx456, nx464, nx520, nx528, nx532, nx544, 
      nx548, nx674, nx678, nx688, nx692, nx756, nx766, nx770, nx776, nx780, 
      nx896, nx900, nx910, nx914, nx978, nx998, nx1002, nx1008, nx1012, 
      nx1118, nx1122, nx1132, nx1136, nx1200, nx1230, nx1234, nx1240, nx1244, 
      nx1340, nx1344, nx1354, nx1358, nx1422, nx1462, nx1466, nx1472, nx1476, 
      nx1562, nx1566, nx1576, nx1580, nx1644, nx1694, nx1698, nx1704, nx1708, 
      nx1784, nx1788, nx1798, nx1802, nx1866, nx1926, nx1930, nx1936, nx1940, 
      nx2006, nx2010, nx2020, nx2024, nx2088, nx2158, nx2162, nx2168, nx2172, 
      nx2228, nx2232, nx2242, nx2246, nx2310, nx2390, nx2394, nx2400, nx2404, 
      nx2450, nx2454, nx2464, nx2468, nx2532, nx2622, nx2626, nx2632, nx2636, 
      nx2672, nx2676, nx2686, nx2690, nx2754, nx2854, nx2858, nx2864, nx2868, 
      nx2894, nx2898, nx2908, nx2912, nx2976, nx3086, nx3090, nx3096, nx3100, 
      nx3116, nx3120, nx3130, nx3134, nx3198, nx3318, nx3322, nx3328, nx3332, 
      nx3338, nx3342, nx3352, nx3356, nx3360, nx3364, nx3420, nx3540, nx3544, 
      nx3574, nx3636, mac_unit_tempP_30, nx1887, mac_unit_tempP_29, nx1889, 
      mac_unit_tempP_28, nx1891, mac_unit_tempP_27, nx1892, 
      mac_unit_tempP_26, nx1893, mac_unit_tempP_25, nx1895, 
      mac_unit_tempP_24, nx1897, mac_unit_tempP_23, nx1899, 
      mac_unit_tempP_22, nx1901, mac_unit_tempP_21, nx1902, 
      mac_unit_tempP_20, nx1903, mac_unit_tempP_19, nx1905, 
      mac_unit_tempP_18, nx1907, mac_unit_tempP_17, nx1909, 
      mac_unit_tempP_16, nx1911, mac_unit_tempP_15, nx1912, 
      mac_unit_tempP_14, nx1913, mac_unit_tempP_13, nx1915, 
      mac_unit_tempP_12, nx1917, mac_unit_tempP_11, nx1919, 
      mac_unit_tempP_10, nx1921, mac_unit_tempP_9, nx1922, mac_unit_tempP_8, 
      nx1923, mac_unit_tempP_7, nx1925, mac_unit_tempP_6, nx1927, 
      mac_unit_tempP_5, nx1929, mac_unit_tempP_4, nx1931, mac_unit_tempP_3, 
      nx1932, mac_unit_tempP_2, nx1933, mac_unit_tempP_1, nx1935, 
      mac_unit_tempP_0, nx1937, nx3638, nx3654, nx3664, nx3678, nx3680, 
      nx3692, nx3702, nx3704, nx3716, nx3726, nx3728, nx3740, nx3750, nx3752, 
      nx3764, nx3774, nx3776, nx3788, nx3798, nx3800, nx3812, nx3822, nx3824, 
      nx3836, nx3846, nx3848, nx3860, nx3870, nx3872, nx3884, nx3894, nx3896, 
      nx3908, nx3918, nx3920, nx3932, nx3942, nx3944, nx3956, nx3966, nx3968, 
      nx3980, nx3990, nx3992, nx4004, nx4014, nx4016, nx4022, nx4034, nx4050, 
      nx4052, nx4058, nx4070, nx4088, nx4106, nx4124, nx4142, nx4160, nx4178, 
      nx4196, nx4214, nx4232, nx4250, nx4268, nx4294, nx4310, nx4318, nx4326, 
      nx4334, nx4342, nx4350, nx4358, nx4366, nx4374, nx4382, nx4390, nx4398, 
      nx4406, nx4414, nx4422, nx4438, sig_0, test_output_misr_signal_31, 
      test_output_misr_signal_30, test_output_misr_signal_29, 
      test_output_misr_signal_28, test_output_misr_signal_27, 
      test_output_misr_signal_26, test_output_misr_signal_25, 
      test_output_misr_signal_24, test_output_misr_signal_23, 
      test_output_misr_signal_22, test_output_misr_signal_21, 
      test_output_misr_signal_20, test_output_misr_signal_19, 
      test_output_misr_signal_18, test_output_misr_signal_17, 
      test_output_misr_signal_16, test_output_misr_signal_15, 
      test_output_misr_signal_14, test_output_misr_signal_13, 
      test_output_misr_signal_12, test_output_misr_signal_11, 
      test_output_misr_signal_10, test_output_misr_signal_9, 
      test_output_misr_signal_8, test_output_misr_signal_7, 
      test_output_misr_signal_6, test_output_misr_signal_5, 
      test_output_misr_signal_4, test_output_misr_signal_3, 
      test_output_misr_signal_2, test_output_misr_signal_1, 
      test_output_misr_signal_0, nx4542, nx4544, nx4550, nx4556, nx4562, 
      nx4568, nx4574, nx4580, nx4586, nx4592, nx4598, nx4604, nx4610, nx4616, 
      nx4628, nx4724, sig_1, sig_2, sig_3, sig_4, sig_5, sig_6, sig_7, sig_8, 
      sig_9, sig_10, sig_11, sig_12, sig_13, sig_14, sig_15, sig_16, sig_17, 
      sig_18, sig_19, sig_20, sig_21, sig_22, sig_23, sig_24, sig_25, sig_26, 
      sig_27, sig_28, sig_29, sig_30, sig_31, nx1945, nx1955, nx1965, nx1975, 
      nx1985, nx1995, nx2005, nx2015, nx2025, nx2035, nx2045, nx2055, nx2065, 
      nx2075, nx2085, nx2095, nx2105, nx2115, nx2125, nx2135, nx2145, nx2155, 
      nx2165, nx2175, nx2185, nx2195, nx2205, nx2215, nx2225, nx2235, nx2245, 
      nx2255, nx2265, nx2275, nx2285, nx2295, nx2305, nx2315, nx2325, nx2335, 
      nx2345, nx2355, nx2365, nx2375, nx2385, nx2395, nx2405, nx2415, nx2429, 
      nx2439, nx2509, nx2513, nx2517, nx2523, nx2555, nx2565, nx2567, nx2579, 
      nx2583, nx2587, nx2591, nx2595, nx2601, nx2603, nx2609, nx2613, nx2621, 
      nx2623, nx2625, nx2627, nx2635, nx2643, nx2645, nx2651, nx2661, nx2668, 
      nx2673, nx2679, nx2681, nx2683, nx2691, nx2699, nx2701, nx2707, nx2717, 
      nx2725, nx2729, nx2735, nx2737, nx2739, nx2741, nx2743, nx2745, nx2747, 
      nx2749, nx2757, nx2765, nx2767, nx2773, nx2783, nx2790, nx2795, nx2801, 
      nx2803, nx2805, nx2807, nx2809, nx2811, nx2813, nx2815, nx2817, nx2819, 
      nx2821, nx2823, nx2831, nx2839, nx2841, nx2847, nx2857, nx2865, nx2869, 
      nx2875, nx2877, nx2879, nx2881, nx2883, nx2885, nx2887, nx2889, nx2891, 
      nx2893, nx2895, nx2897, nx2899, nx2901, nx2903, nx2905, nx2913, nx2921, 
      nx2923, nx2929, nx2939, nx2947, nx2951, nx2957, nx2959, nx2961, nx2963, 
      nx2965, nx2967, nx2969, nx2971, nx2973, nx2975, nx2977, nx2979, nx2981, 
      nx2983, nx2985, nx2987, nx2989, nx2991, nx2993, nx2995, nx3003, nx3011, 
      nx3013, nx3019, nx3029, nx3033, nx3037, nx3043, nx3045, nx3047, nx3049, 
      nx3051, nx3053, nx3055, nx3057, nx3059, nx3061, nx3063, nx3065, nx3067, 
      nx3069, nx3071, nx3073, nx3075, nx3077, nx3079, nx3081, nx3083, nx3085, 
      nx3087, nx3089, nx3095, nx3103, nx3105, nx3111, nx3121, nx3125, nx3129, 
      nx3135, nx3137, nx3139, nx3141, nx3143, nx3145, nx3147, nx3149, nx3151, 
      nx3153, nx3155, nx3157, nx3159, nx3161, nx3163, nx3165, nx3167, nx3169, 
      nx3171, nx3173, nx3175, nx3177, nx3179, nx3181, nx3183, nx3185, nx3187, 
      nx3189, nx3195, nx3203, nx3205, nx3211, nx3221, nx3225, nx3229, nx3235, 
      nx3237, nx3239, nx3241, nx3243, nx3245, nx3247, nx3249, nx3251, nx3253, 
      nx3255, nx3257, nx3259, nx3261, nx3263, nx3265, nx3267, nx3269, nx3271, 
      nx3273, nx3275, nx3277, nx3279, nx3281, nx3283, nx3285, nx3287, nx3289, 
      nx3291, nx3293, nx3295, nx3297, nx3303, nx3311, nx3313, nx3319, nx3329, 
      nx3333, nx3337, nx3343, nx3345, nx3347, nx3349, nx3351, nx3353, nx3355, 
      nx3357, nx3359, nx3361, nx3363, nx3365, nx3367, nx3369, nx3371, nx3373, 
      nx3375, nx3377, nx3379, nx3381, nx3383, nx3385, nx3387, nx3389, nx3391, 
      nx3393, nx3395, nx3397, nx3399, nx3401, nx3403, nx3405, nx3407, nx3409, 
      nx3411, nx3413, nx3417, nx3425, nx3427, nx3433, nx3443, nx3447, nx3451, 
      nx3457, nx3459, nx3461, nx3463, nx3465, nx3467, nx3469, nx3471, nx3473, 
      nx3475, nx3477, nx3479, nx3481, nx3483, nx3485, nx3487, nx3489, nx3491, 
      nx3493, nx3495, nx3497, nx3499, nx3501, nx3503, nx3505, nx3507, nx3509, 
      nx3511, nx3513, nx3515, nx3517, nx3519, nx3521, nx3523, nx3525, nx3527, 
      nx3529, nx3531, nx3533, nx3535, nx3541, nx3549, nx3551, nx3557, nx3567, 
      nx3571, nx3575, nx3581, nx3583, nx3585, nx3587, nx3589, nx3591, nx3593, 
      nx3595, nx3597, nx3599, nx3601, nx3603, nx3605, nx3607, nx3609, nx3611, 
      nx3613, nx3615, nx3617, nx3619, nx3621, nx3623, nx3625, nx3627, nx3629, 
      nx3631, nx3633, nx3635, nx3637, nx3639, nx3641, nx3643, nx3645, nx3647, 
      nx3649, nx3651, nx3653, nx3655, nx3657, nx3659, nx3661, nx3663, nx3665, 
      nx3667, nx3673, nx3681, nx3683, nx3687, nx3697, nx3701, nx3705, nx3709, 
      nx3711, nx3713, nx3715, nx3717, nx3719, nx3721, nx3723, nx3725, nx3727, 
      nx3729, nx3731, nx3733, nx3735, nx3737, nx3739, nx3741, nx3743, nx3745, 
      nx3747, nx3749, nx3751, nx3753, nx3755, nx3757, nx3759, nx3761, nx3763, 
      nx3765, nx3767, nx3769, nx3771, nx3773, nx3775, nx3777, nx3779, nx3781, 
      nx3783, nx3785, nx3787, nx3789, nx3791, nx3793, nx3795, nx3797, nx3799, 
      nx3801, nx3803, nx3807, nx3815, nx3817, nx3823, nx3833, nx3837, nx3841, 
      nx3847, nx3849, nx3851, nx3853, nx3855, nx3857, nx3859, nx3861, nx3863, 
      nx3865, nx3867, nx3869, nx3871, nx3873, nx3875, nx3877, nx3879, nx3881, 
      nx3883, nx3885, nx3887, nx3889, nx3891, nx3893, nx3895, nx3897, nx3899, 
      nx3901, nx3903, nx3905, nx3907, nx3909, nx3911, nx3913, nx3915, nx3917, 
      nx3919, nx3921, nx3923, nx3925, nx3927, nx3929, nx3931, nx3933, nx3935, 
      nx3937, nx3939, nx3941, nx3943, nx3945, nx3947, nx3949, nx3955, nx3963, 
      nx3965, nx3971, nx3979, nx3981, nx3983, nx3989, nx3993, nx3995, nx3999, 
      nx4003, nx4007, nx4011, nx4015, nx4019, nx4023, nx4027, nx4031, nx4035, 
      nx4038, nx4041, nx4045, nx4049, nx4053, nx4056, nx4059, nx4063, nx4067, 
      nx4071, nx4074, nx4077, nx4081, nx4085, nx4087, nx4091, nx4095, nx4105, 
      nx4107, nx4109, nx4111, nx4113, nx4115, nx4121, nx4125, nx4127, nx4131, 
      nx4135, nx4137, nx4141, nx4145, nx4147, nx4151, nx4155, nx4157, nx4161, 
      nx4164, nx4167, nx4171, nx4175, nx4177, nx4181, nx4185, nx4187, nx4191, 
      nx4195, nx4197, nx4200, nx4203, nx4205, nx4209, nx4213, nx4215, nx4218, 
      nx4221, nx4223, nx4227, nx4231, nx4233, nx4237, nx4239, nx4251, nx4253, 
      nx4257, nx4261, nx4265, nx4271, nx4273, nx4275, nx4277, nx4279, nx4281, 
      nx4283, nx4285, nx4287, nx4289, nx4291, nx4293, nx4295, nx4297, nx4299, 
      nx4301, nx4303, nx4305, nx4307, nx4309, nx4311, nx4313, nx4315, nx4317, 
      nx4319, nx4321, nx4323, nx4325, nx4327, nx4329, nx4331, nx4333, nx4335, 
      nx4337, nx4339, nx4341, nx4343, nx4345, nx4347, nx4349, nx4351, nx4353, 
      nx4355, nx4357, nx4359, nx4361, nx4363, nx4365, nx4367, nx4369, nx4371, 
      nx4373, nx4375, nx4377, nx4379, nx4381, nx4383, nx4385, nx4387, nx4391, 
      nx4399, nx4401, nx4403, nx4405, nx4407, nx4409, nx4411, nx4413, nx4415, 
      nx4417, nx4419, nx4421, nx4423, nx4425, nx4427, nx4429, nx4431, nx4433, 
      nx4435, nx4437, nx4439, nx4441, nx4443, nx4445, nx4447, nx4449, nx4451, 
      nx4453, nx4455, nx4457, nx4459, nx4461, nx4463, nx4465, nx4467, nx4469, 
      nx4471, nx4473, nx4475, nx4477, nx4479, nx4481, nx4483, nx4485, nx4487, 
      nx4489, nx4491, nx4493, nx4495, nx4497, nx4499, nx4501, nx4511, nx4519, 
      nx4521, nx4523, nx4525, nx4527, nx4529, nx4531, nx4533, nx4535, nx4537, 
      nx4539, nx4541, nx4543, nx4545, nx4547, nx4549, nx4551, nx4553, nx4555, 
      nx4557, nx4559, nx4561, nx4563, nx4565, nx4567, nx4569, nx4571, nx4573, 
      nx4575, nx4577, nx4579, nx4581, nx4583, nx4585, nx4587, nx4589, nx4591, 
      nx4593, nx4595, nx4597, nx4599, nx4601, nx4603, nx4605, nx4607, nx4609, 
      nx4613, nx4620, nx4623, nx4625, nx4627, nx4629, nx4631, nx4633, nx4635, 
      nx4637, nx4639, nx4641, nx4643, nx4645, nx4647, nx4649, nx4651, nx4653, 
      nx4655, nx4657, nx4659, nx4661, nx4663, nx4665, nx4667, nx4669, nx4671, 
      nx4673, nx4675, nx4677, nx4679, nx4681, nx4683, nx4685, nx4687, nx4689, 
      nx4691, nx4693, nx4695, nx4697, nx4699, nx4701, nx4703, nx4707, nx4714, 
      nx4716, nx4719, nx4721, nx4723, nx4725, nx4727, nx4729, nx4731, nx4733, 
      nx4735, nx4737, nx4739, nx4741, nx4743, nx4745, nx4747, nx4749, nx4751, 
      nx4753, nx4755, nx4757, nx4759, nx4761, nx4763, nx4765, nx4767, nx4769, 
      nx4771, nx4773, nx4775, nx4777, nx4779, nx4781, nx4783, nx4785, nx4787, 
      nx4789, nx4793, nx4799, nx4801, nx4803, nx4805, nx4807, nx4809, nx4811, 
      nx4813, nx4815, nx4817, nx4819, nx4821, nx4823, nx4825, nx4827, nx4829, 
      nx4831, nx4833, nx4835, nx4837, nx4839, nx4841, nx4843, nx4845, nx4847, 
      nx4849, nx4851, nx4853, nx4855, nx4857, nx4859, nx4861, nx4863, nx4865, 
      nx4868, nx4875, nx4877, nx4879, nx4881, nx4883, nx4885, nx4887, nx4889, 
      nx4891, nx4893, nx4895, nx4897, nx4899, nx4901, nx4903, nx4905, nx4907, 
      nx4909, nx4911, nx4913, nx4915, nx4917, nx4919, nx4921, nx4923, nx4925, 
      nx4927, nx4929, nx4931, nx4933, nx4937, nx4943, nx4945, nx4947, nx4949, 
      nx4951, nx4953, nx4955, nx4957, nx4959, nx4961, nx4963, nx4965, nx4967, 
      nx4969, nx4971, nx4973, nx4975, nx4977, nx4979, nx4981, nx4983, nx4985, 
      nx4987, nx4989, nx4991, nx4993, nx4996, nx5002, nx5004, nx5006, nx5008, 
      nx5010, nx5012, nx5014, nx5016, nx5018, nx5020, nx5022, nx5024, nx5026, 
      nx5028, nx5030, nx5032, nx5034, nx5036, nx5038, nx5040, nx5042, nx5044, 
      nx5047, nx5053, nx5055, nx5057, nx5059, nx5061, nx5063, nx5065, nx5067, 
      nx5069, nx5071, nx5073, nx5075, nx5077, nx5079, nx5081, nx5083, nx5085, 
      nx5087, nx5090, nx5096, nx5098, nx5100, nx5102, nx5104, nx5106, nx5108, 
      nx5110, nx5112, nx5114, nx5116, nx5118, nx5120, nx5122, nx5125, nx5131, 
      nx5133, nx5135, nx5137, nx5139, nx5141, nx5143, nx5145, nx5147, nx5149, 
      nx5152, nx5158, nx5160, nx5162, nx5164, nx5166, nx5168, nx5175, nx5177, 
      nx5183, nx5191, nx5195, nx5199, nx5203, nx5207, nx5211, nx5215, nx5219, 
      nx5223, nx5227, nx5231, nx5235, nx5239, nx5243, nx5247, nx5254, nx5296, 
      nx5311, nx5314, nx5316, nx5318, nx5320, nx5322, nx5324, nx5326, nx5328, 
      nx5330, nx5332, nx5334, nx5336, nx5338, nx5340, nx5342, nx5345, nx5446, 
      nx5448, nx5450, nx5456, nx5464, nx5468, nx5472, nx5476, nx5480, nx5484, 
      nx5488, nx5492, nx5496, nx5500, nx5504, nx5508, nx5512, nx5516, nx5520, 
      nx5524, nx5526, nx5534, nx5536, nx5542, nx5544, nx5546, nx5548, nx5550
   : std_logic ;

begin
   ix4299 : nor02 port map ( Y=>mac_output(0), A0=>RST, A1=>nx2429);
   ix2430 : xnor2 port map ( Y=>nx2429, A0=>Cin, A1=>nx1937);
   ix3645 : xnor2 port map ( Y=>nx1937, A0=>mac_unit_tempP_0, A1=>nx2439);
   mac_unit_MR_reg_Q_0 : dffr port map ( Q=>mac_unit_tempP_0, QB=>OPEN, D=>
      nx3638, CLK=>CLK, R=>RST);
   ix91 : mux21 port map ( Y=>nx90, A0=>B(0), A1=>lfsr_C_15, S0=>test_mode);
   test_input_reg_BP2_15 : dff port map ( Q=>lfsr_C_15, QB=>OPEN, D=>
      test_input_lfsr_signal_15, CLK=>CLK);
   test_input_reg_lfsr_signal_15 : dffs port map ( Q=>
      test_input_lfsr_signal_15, QB=>OPEN, D=>nx2095, CLK=>CLK, S=>RST);
   test_input_reg_lfsr_signal_14 : dffr port map ( Q=>
      test_input_lfsr_signal_14, QB=>OPEN, D=>nx2085, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_13 : dffr port map ( Q=>
      test_input_lfsr_signal_13, QB=>OPEN, D=>nx2075, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_12 : dffr port map ( Q=>
      test_input_lfsr_signal_12, QB=>OPEN, D=>nx2065, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_11 : dffr port map ( Q=>
      test_input_lfsr_signal_11, QB=>OPEN, D=>nx2055, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_10 : dffr port map ( Q=>
      test_input_lfsr_signal_10, QB=>OPEN, D=>nx2045, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_9 : dffr port map ( Q=>
      test_input_lfsr_signal_9, QB=>OPEN, D=>nx2035, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_8 : dffr port map ( Q=>
      test_input_lfsr_signal_8, QB=>OPEN, D=>nx2025, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_7 : dffr port map ( Q=>
      test_input_lfsr_signal_7, QB=>OPEN, D=>nx2015, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_6 : dffr port map ( Q=>
      test_input_lfsr_signal_6, QB=>OPEN, D=>nx2005, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_5 : dffr port map ( Q=>
      test_input_lfsr_signal_5, QB=>OPEN, D=>nx1995, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_4 : dffr port map ( Q=>
      test_input_lfsr_signal_4, QB=>OPEN, D=>nx1985, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_3 : dffr port map ( Q=>
      test_input_lfsr_signal_3, QB=>OPEN, D=>nx1975, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_2 : dffr port map ( Q=>
      test_input_lfsr_signal_2, QB=>OPEN, D=>nx1965, CLK=>CLK, R=>RST);
   test_input_reg_lfsr_signal_1 : dffr port map ( Q=>
      test_input_lfsr_signal_1, QB=>OPEN, D=>nx1955, CLK=>CLK, R=>RST);
   ix1946 : oai32 port map ( Y=>nx1945, A0=>nx2509, A1=>RST, A2=>nx5524, B0
      =>nx2517, B1=>nx5446);
   ix2510 : xnor2 port map ( Y=>nx2509, A0=>test_input_lfsr_signal_10, A1=>
      nx14);
   ix15 : xnor2 port map ( Y=>nx14, A0=>test_input_lfsr_signal_12, A1=>
      nx2513);
   ix2514 : xnor2 port map ( Y=>nx2513, A0=>test_input_lfsr_signal_15, A1=>
      test_input_lfsr_signal_13);
   test_input_reg_lfsr_signal_0 : dffr port map ( Q=>
      test_input_lfsr_signal_0, QB=>nx2517, D=>nx1945, CLK=>CLK, R=>RST);
   ix2524 : inv01 port map ( Y=>nx2523, A=>RST);
   ix457 : mux21 port map ( Y=>nx456, A0=>C(0), A1=>lfsr_B_15, S0=>test_mode
   );
   test_input_reg_BP1_15 : dff port map ( Q=>lfsr_B_15, QB=>OPEN, D=>
      test_input_lfsr_signal_0, CLK=>CLK);
   ix4307 : nor02 port map ( Y=>mac_output(1), A0=>RST, A1=>nx2555);
   ix2556 : nand02 port map ( Y=>nx2555, A0=>nx2523, A1=>nx3654);
   ix3655 : xnor2 port map ( Y=>nx3654, A0=>nx1935, A1=>nx2595);
   ix3671 : xnor2 port map ( Y=>nx1935, A0=>mac_unit_tempP_1, A1=>nx2565);
   mac_unit_MR_reg_Q_1 : dffr port map ( Q=>mac_unit_tempP_1, QB=>OPEN, D=>
      nx3654, CLK=>CLK, R=>RST);
   ix2566 : nand02 port map ( Y=>nx2565, A0=>nx2567, A1=>nx3664);
   ix115 : mux21 port map ( Y=>nx114, A0=>B(1), A1=>lfsr_C_14, S0=>test_mode
   );
   test_input_reg_BP2_14 : dff port map ( Q=>lfsr_C_14, QB=>OPEN, D=>
      test_input_lfsr_signal_14, CLK=>CLK);
   ix435 : mux21 port map ( Y=>nx434, A0=>C(1), A1=>lfsr_C_1, S0=>test_mode
   );
   test_input_reg_BP2_1 : dff port map ( Q=>lfsr_C_1, QB=>OPEN, D=>
      test_input_lfsr_signal_1, CLK=>CLK);
   ix2596 : aoi32 port map ( Y=>nx2595, A0=>nx5448, A1=>nx5464, A2=>
      mac_unit_tempP_0, B0=>Cin, B1=>nx1937);
   ix4315 : nor02ii port map ( Y=>mac_output(2), A0=>RST, A1=>nx4310);
   ix4311 : nor02 port map ( Y=>nx4310, A0=>RST, A1=>nx2601);
   ix2602 : xnor2 port map ( Y=>nx2601, A0=>nx2603, A1=>nx2609);
   ix2604 : xnor2 port map ( Y=>nx2603, A0=>mac_unit_tempP_2, A1=>nx3692);
   mac_unit_MR_reg_Q_2 : dffr port map ( Q=>mac_unit_tempP_2, QB=>OPEN, D=>
      nx3680, CLK=>CLK, R=>RST);
   ix2610 : mux21 port map ( Y=>nx2609, A0=>nx2565, A1=>nx2595, S0=>nx1935);
   ix3693 : aoi21 port map ( Y=>nx3692, A0=>nx2613, A1=>nx2621, B0=>nx688);
   ix529 : mux21 port map ( Y=>nx528, A0=>B(2), A1=>lfsr_C_13, S0=>test_mode
   );
   test_input_reg_BP2_13 : dff port map ( Q=>lfsr_C_13, QB=>OPEN, D=>
      test_input_lfsr_signal_13, CLK=>CLK);
   ix2622 : xnor2 port map ( Y=>nx2621, A0=>nx2567, A1=>nx2623);
   ix2624 : xnor2 port map ( Y=>nx2623, A0=>nx2625, A1=>nx2627);
   ix2628 : nand02 port map ( Y=>nx2627, A0=>nx5448, A1=>nx410);
   ix411 : mux21 port map ( Y=>nx410, A0=>C(2), A1=>lfsr_C_2, S0=>test_mode
   );
   test_input_reg_BP2_2 : dff port map ( Q=>lfsr_C_2, QB=>OPEN, D=>
      test_input_lfsr_signal_2, CLK=>CLK);
   ix689 : nor03 port map ( Y=>nx688, A0=>nx2621, A1=>nx5536, A2=>nx2635);
   ix4323 : nor02ii port map ( Y=>mac_output(3), A0=>RST, A1=>nx4318);
   ix4319 : nor02 port map ( Y=>nx4318, A0=>RST, A1=>nx2643);
   ix2644 : xnor2 port map ( Y=>nx2643, A0=>nx2645, A1=>nx2651);
   ix2646 : xnor2 port map ( Y=>nx2645, A0=>mac_unit_tempP_3, A1=>nx3716);
   mac_unit_MR_reg_Q_3 : dffr port map ( Q=>mac_unit_tempP_3, QB=>OPEN, D=>
      nx3704, CLK=>CLK, R=>RST);
   ix2652 : aoi22 port map ( Y=>nx2651, A0=>nx3692, A1=>mac_unit_tempP_2, B0
      =>nx1933, B1=>nx3678);
   ix3717 : aoi21 port map ( Y=>nx3716, A0=>nx2661, A1=>nx2668, B0=>nx910);
   ix757 : mux21 port map ( Y=>nx756, A0=>B(3), A1=>lfsr_C_12, S0=>test_mode
   );
   test_input_reg_BP2_12 : dff port map ( Q=>lfsr_C_12, QB=>OPEN, D=>
      test_input_lfsr_signal_12, CLK=>CLK);
   ix2670 : xnor2 port map ( Y=>nx2668, A0=>nx688, A1=>nx678);
   ix679 : xnor2 port map ( Y=>nx678, A0=>nx2673, A1=>nx674);
   ix675 : xnor2 port map ( Y=>nx674, A0=>nx464, A1=>nx2679);
   ix465 : aoi21 port map ( Y=>nx464, A0=>nx2439, A1=>nx2627, B0=>nx2625);
   ix2680 : xnor2 port map ( Y=>nx2679, A0=>nx2681, A1=>nx2683);
   ix2682 : nand02 port map ( Y=>nx2681, A0=>nx5456, A1=>nx410);
   ix2684 : nand02 port map ( Y=>nx2683, A0=>nx5448, A1=>nx386);
   ix387 : mux21 port map ( Y=>nx386, A0=>C(3), A1=>lfsr_C_3, S0=>test_mode
   );
   test_input_reg_BP2_3 : dff port map ( Q=>lfsr_C_3, QB=>OPEN, D=>
      test_input_lfsr_signal_3, CLK=>CLK);
   ix911 : nor03 port map ( Y=>nx910, A0=>nx2668, A1=>nx5536, A2=>nx2691);
   ix4331 : nor02ii port map ( Y=>mac_output(4), A0=>RST, A1=>nx4326);
   ix4327 : nor02 port map ( Y=>nx4326, A0=>RST, A1=>nx2699);
   ix2700 : xnor2 port map ( Y=>nx2699, A0=>nx2701, A1=>nx2707);
   ix2702 : xnor2 port map ( Y=>nx2701, A0=>mac_unit_tempP_4, A1=>nx3740);
   mac_unit_MR_reg_Q_4 : dffr port map ( Q=>mac_unit_tempP_4, QB=>OPEN, D=>
      nx3728, CLK=>CLK, R=>RST);
   ix2708 : aoi22 port map ( Y=>nx2707, A0=>nx3716, A1=>mac_unit_tempP_3, B0
      =>nx1932, B1=>nx3702);
   ix3741 : aoi21 port map ( Y=>nx3740, A0=>nx2717, A1=>nx2725, B0=>nx1132);
   ix979 : mux21 port map ( Y=>nx978, A0=>B(4), A1=>lfsr_C_11, S0=>test_mode
   );
   test_input_reg_BP2_11 : dff port map ( Q=>lfsr_C_11, QB=>OPEN, D=>
      test_input_lfsr_signal_11, CLK=>CLK);
   ix2726 : xnor2 port map ( Y=>nx2725, A0=>nx910, A1=>nx900);
   ix901 : xnor2 port map ( Y=>nx900, A0=>nx2729, A1=>nx896);
   ix897 : xnor2 port map ( Y=>nx896, A0=>nx692, A1=>nx2735);
   ix693 : mux21 port map ( Y=>nx692, A0=>nx674, A1=>nx688, S0=>nx678);
   ix2736 : xnor2 port map ( Y=>nx2735, A0=>nx2737, A1=>nx2739);
   ix2738 : nand02 port map ( Y=>nx2737, A0=>nx5468, A1=>nx410);
   ix2740 : xnor2 port map ( Y=>nx2739, A0=>nx2741, A1=>nx2745);
   ix2742 : mux21 port map ( Y=>nx2741, A0=>nx2743, A1=>nx2683, S0=>nx2679);
   ix2746 : xnor2 port map ( Y=>nx2745, A0=>nx2747, A1=>nx2749);
   ix2748 : nand02 port map ( Y=>nx2747, A0=>nx5456, A1=>nx386);
   ix2750 : nand02 port map ( Y=>nx2749, A0=>nx5448, A1=>nx362);
   ix363 : mux21 port map ( Y=>nx362, A0=>C(4), A1=>lfsr_C_4, S0=>test_mode
   );
   test_input_reg_BP2_4 : dff port map ( Q=>lfsr_C_4, QB=>OPEN, D=>
      test_input_lfsr_signal_4, CLK=>CLK);
   ix1133 : nor03 port map ( Y=>nx1132, A0=>nx2725, A1=>nx5536, A2=>nx2757);
   ix4339 : nor02ii port map ( Y=>mac_output(5), A0=>RST, A1=>nx4334);
   ix4335 : nor02 port map ( Y=>nx4334, A0=>RST, A1=>nx2765);
   ix2766 : xnor2 port map ( Y=>nx2765, A0=>nx2767, A1=>nx2773);
   ix2768 : xnor2 port map ( Y=>nx2767, A0=>mac_unit_tempP_5, A1=>nx3764);
   mac_unit_MR_reg_Q_5 : dffr port map ( Q=>mac_unit_tempP_5, QB=>OPEN, D=>
      nx3752, CLK=>CLK, R=>RST);
   ix2774 : aoi22 port map ( Y=>nx2773, A0=>nx3740, A1=>mac_unit_tempP_4, B0
      =>nx1931, B1=>nx3726);
   ix3765 : aoi21 port map ( Y=>nx3764, A0=>nx2783, A1=>nx2790, B0=>nx1354);
   ix1201 : mux21 port map ( Y=>nx1200, A0=>B(5), A1=>lfsr_C_10, S0=>
      test_mode);
   test_input_reg_BP2_10 : dff port map ( Q=>lfsr_C_10, QB=>OPEN, D=>
      test_input_lfsr_signal_10, CLK=>CLK);
   ix2792 : xnor2 port map ( Y=>nx2790, A0=>nx1132, A1=>nx1122);
   ix1123 : xnor2 port map ( Y=>nx1122, A0=>nx2795, A1=>nx1118);
   ix1119 : xnor2 port map ( Y=>nx1118, A0=>nx914, A1=>nx2801);
   ix915 : mux21 port map ( Y=>nx914, A0=>nx896, A1=>nx910, S0=>nx900);
   ix2802 : xnor2 port map ( Y=>nx2801, A0=>nx2803, A1=>nx2805);
   ix2804 : nand02 port map ( Y=>nx2803, A0=>nx410, A1=>nx5472);
   ix2806 : xnor2 port map ( Y=>nx2805, A0=>nx2807, A1=>nx2811);
   ix2808 : mux21 port map ( Y=>nx2807, A0=>nx2809, A1=>nx2739, S0=>nx2735);
   ix2812 : xnor2 port map ( Y=>nx2811, A0=>nx2813, A1=>nx2815);
   ix2814 : nand02 port map ( Y=>nx2813, A0=>nx5468, A1=>nx386);
   ix2816 : xnor2 port map ( Y=>nx2815, A0=>nx2817, A1=>nx2819);
   ix2818 : mux21 port map ( Y=>nx2817, A0=>nx2741, A1=>nx2749, S0=>nx2745);
   ix2820 : xnor2 port map ( Y=>nx2819, A0=>nx2821, A1=>nx2823);
   ix2822 : nand02 port map ( Y=>nx2821, A0=>nx5456, A1=>nx362);
   ix2824 : nand02 port map ( Y=>nx2823, A0=>nx5448, A1=>nx338);
   ix339 : mux21 port map ( Y=>nx338, A0=>C(5), A1=>lfsr_C_5, S0=>test_mode
   );
   test_input_reg_BP2_5 : dff port map ( Q=>lfsr_C_5, QB=>OPEN, D=>
      test_input_lfsr_signal_5, CLK=>CLK);
   ix1355 : nor03 port map ( Y=>nx1354, A0=>nx2790, A1=>nx5536, A2=>nx2831);
   ix4347 : nor02ii port map ( Y=>mac_output(6), A0=>RST, A1=>nx4342);
   ix4343 : nor02 port map ( Y=>nx4342, A0=>RST, A1=>nx2839);
   ix2840 : xnor2 port map ( Y=>nx2839, A0=>nx2841, A1=>nx2847);
   ix2842 : xnor2 port map ( Y=>nx2841, A0=>mac_unit_tempP_6, A1=>nx3788);
   mac_unit_MR_reg_Q_6 : dffr port map ( Q=>mac_unit_tempP_6, QB=>OPEN, D=>
      nx3776, CLK=>CLK, R=>RST);
   ix2848 : aoi22 port map ( Y=>nx2847, A0=>nx3764, A1=>mac_unit_tempP_5, B0
      =>nx1929, B1=>nx3750);
   ix3789 : aoi21 port map ( Y=>nx3788, A0=>nx2857, A1=>nx2865, B0=>nx1576);
   ix1423 : mux21 port map ( Y=>nx1422, A0=>B(6), A1=>lfsr_C_9, S0=>
      test_mode);
   test_input_reg_BP2_9 : dff port map ( Q=>lfsr_C_9, QB=>OPEN, D=>
      test_input_lfsr_signal_9, CLK=>CLK);
   ix2866 : xnor2 port map ( Y=>nx2865, A0=>nx1354, A1=>nx1344);
   ix1345 : xnor2 port map ( Y=>nx1344, A0=>nx2869, A1=>nx1340);
   ix1341 : xnor2 port map ( Y=>nx1340, A0=>nx1136, A1=>nx2875);
   ix1137 : mux21 port map ( Y=>nx1136, A0=>nx1118, A1=>nx1132, S0=>nx1122);
   ix2876 : xnor2 port map ( Y=>nx2875, A0=>nx2877, A1=>nx2879);
   ix2878 : nand02 port map ( Y=>nx2877, A0=>nx410, A1=>nx5476);
   ix2880 : xnor2 port map ( Y=>nx2879, A0=>nx2881, A1=>nx2885);
   ix2882 : mux21 port map ( Y=>nx2881, A0=>nx2883, A1=>nx2805, S0=>nx2801);
   ix2886 : xnor2 port map ( Y=>nx2885, A0=>nx2887, A1=>nx2889);
   ix2888 : nand02 port map ( Y=>nx2887, A0=>nx5472, A1=>nx386);
   ix2890 : xnor2 port map ( Y=>nx2889, A0=>nx2891, A1=>nx2893);
   ix2892 : mux21 port map ( Y=>nx2891, A0=>nx2807, A1=>nx2815, S0=>nx2811);
   ix2894 : xnor2 port map ( Y=>nx2893, A0=>nx2895, A1=>nx2897);
   ix2896 : nand02 port map ( Y=>nx2895, A0=>nx5468, A1=>nx362);
   ix2898 : xnor2 port map ( Y=>nx2897, A0=>nx2899, A1=>nx2901);
   ix2900 : mux21 port map ( Y=>nx2899, A0=>nx2817, A1=>nx2823, S0=>nx2819);
   ix2902 : xnor2 port map ( Y=>nx2901, A0=>nx2903, A1=>nx2905);
   ix2904 : nand02 port map ( Y=>nx2903, A0=>nx5456, A1=>nx338);
   ix2906 : nand02 port map ( Y=>nx2905, A0=>nx5448, A1=>nx314);
   ix315 : mux21 port map ( Y=>nx314, A0=>C(6), A1=>lfsr_C_6, S0=>test_mode
   );
   test_input_reg_BP2_6 : dff port map ( Q=>lfsr_C_6, QB=>OPEN, D=>
      test_input_lfsr_signal_6, CLK=>CLK);
   ix1577 : nor03 port map ( Y=>nx1576, A0=>nx2865, A1=>nx5536, A2=>nx2913);
   ix4355 : nor02ii port map ( Y=>mac_output(7), A0=>RST, A1=>nx4350);
   ix4351 : nor02 port map ( Y=>nx4350, A0=>RST, A1=>nx2921);
   ix2922 : xnor2 port map ( Y=>nx2921, A0=>nx2923, A1=>nx2929);
   ix2924 : xnor2 port map ( Y=>nx2923, A0=>mac_unit_tempP_7, A1=>nx3812);
   mac_unit_MR_reg_Q_7 : dffr port map ( Q=>mac_unit_tempP_7, QB=>OPEN, D=>
      nx3800, CLK=>CLK, R=>RST);
   ix2930 : aoi22 port map ( Y=>nx2929, A0=>nx3788, A1=>mac_unit_tempP_6, B0
      =>nx1927, B1=>nx3774);
   ix3813 : aoi21 port map ( Y=>nx3812, A0=>nx2939, A1=>nx2947, B0=>nx1798);
   ix1645 : mux21 port map ( Y=>nx1644, A0=>B(7), A1=>lfsr_C_8, S0=>
      test_mode);
   test_input_reg_BP2_8 : dff port map ( Q=>lfsr_C_8, QB=>OPEN, D=>
      test_input_lfsr_signal_8, CLK=>CLK);
   ix2948 : xnor2 port map ( Y=>nx2947, A0=>nx1576, A1=>nx1566);
   ix1567 : xnor2 port map ( Y=>nx1566, A0=>nx2951, A1=>nx1562);
   ix1563 : xnor2 port map ( Y=>nx1562, A0=>nx1358, A1=>nx2957);
   ix1359 : mux21 port map ( Y=>nx1358, A0=>nx1340, A1=>nx1354, S0=>nx1344);
   ix2958 : xnor2 port map ( Y=>nx2957, A0=>nx2959, A1=>nx2961);
   ix2960 : nand02 port map ( Y=>nx2959, A0=>nx410, A1=>nx5480);
   ix2962 : xnor2 port map ( Y=>nx2961, A0=>nx2963, A1=>nx2967);
   ix2964 : mux21 port map ( Y=>nx2963, A0=>nx2965, A1=>nx2879, S0=>nx2875);
   ix2968 : xnor2 port map ( Y=>nx2967, A0=>nx2969, A1=>nx2971);
   ix2970 : nand02 port map ( Y=>nx2969, A0=>nx386, A1=>nx5476);
   ix2972 : xnor2 port map ( Y=>nx2971, A0=>nx2973, A1=>nx2975);
   ix2974 : mux21 port map ( Y=>nx2973, A0=>nx2881, A1=>nx2889, S0=>nx2885);
   ix2976 : xnor2 port map ( Y=>nx2975, A0=>nx2977, A1=>nx2979);
   ix2978 : nand02 port map ( Y=>nx2977, A0=>nx5472, A1=>nx362);
   ix2980 : xnor2 port map ( Y=>nx2979, A0=>nx2981, A1=>nx2983);
   ix2982 : mux21 port map ( Y=>nx2981, A0=>nx2891, A1=>nx2897, S0=>nx2893);
   ix2984 : xnor2 port map ( Y=>nx2983, A0=>nx2985, A1=>nx2987);
   ix2986 : nand02 port map ( Y=>nx2985, A0=>nx5468, A1=>nx338);
   ix2988 : xnor2 port map ( Y=>nx2987, A0=>nx2989, A1=>nx2991);
   ix2990 : mux21 port map ( Y=>nx2989, A0=>nx2899, A1=>nx2905, S0=>nx2901);
   ix2992 : xnor2 port map ( Y=>nx2991, A0=>nx2993, A1=>nx2995);
   ix2994 : nand02 port map ( Y=>nx2993, A0=>nx5456, A1=>nx314);
   ix2996 : nand02 port map ( Y=>nx2995, A0=>nx5448, A1=>nx290);
   ix291 : mux21 port map ( Y=>nx290, A0=>C(7), A1=>lfsr_C_7, S0=>test_mode
   );
   test_input_reg_BP2_7 : dff port map ( Q=>lfsr_C_7, QB=>OPEN, D=>
      test_input_lfsr_signal_7, CLK=>CLK);
   ix1799 : nor03 port map ( Y=>nx1798, A0=>nx2947, A1=>nx5536, A2=>nx3003);
   ix4363 : nor02ii port map ( Y=>mac_output(8), A0=>RST, A1=>nx4358);
   ix4359 : nor02 port map ( Y=>nx4358, A0=>RST, A1=>nx3011);
   ix3012 : xnor2 port map ( Y=>nx3011, A0=>nx3013, A1=>nx3019);
   ix3014 : xnor2 port map ( Y=>nx3013, A0=>mac_unit_tempP_8, A1=>nx3836);
   mac_unit_MR_reg_Q_8 : dffr port map ( Q=>mac_unit_tempP_8, QB=>OPEN, D=>
      nx3824, CLK=>CLK, R=>RST);
   ix3020 : aoi22 port map ( Y=>nx3019, A0=>nx3812, A1=>mac_unit_tempP_7, B0
      =>nx1925, B1=>nx3798);
   ix3837 : aoi21 port map ( Y=>nx3836, A0=>nx3029, A1=>nx3033, B0=>nx2020);
   ix1867 : mux21 port map ( Y=>nx1866, A0=>B(8), A1=>lfsr_C_7, S0=>
      test_mode);
   ix3034 : xnor2 port map ( Y=>nx3033, A0=>nx1798, A1=>nx1788);
   ix1789 : xnor2 port map ( Y=>nx1788, A0=>nx3037, A1=>nx1784);
   ix1785 : xnor2 port map ( Y=>nx1784, A0=>nx1580, A1=>nx3043);
   ix1581 : mux21 port map ( Y=>nx1580, A0=>nx1562, A1=>nx1576, S0=>nx1566);
   ix3044 : xnor2 port map ( Y=>nx3043, A0=>nx3045, A1=>nx3047);
   ix3046 : nand02 port map ( Y=>nx3045, A0=>nx410, A1=>nx5484);
   ix3048 : xnor2 port map ( Y=>nx3047, A0=>nx3049, A1=>nx3053);
   ix3050 : mux21 port map ( Y=>nx3049, A0=>nx3051, A1=>nx2961, S0=>nx2957);
   ix3054 : xnor2 port map ( Y=>nx3053, A0=>nx3055, A1=>nx3057);
   ix3056 : nand02 port map ( Y=>nx3055, A0=>nx386, A1=>nx5480);
   ix3058 : xnor2 port map ( Y=>nx3057, A0=>nx3059, A1=>nx3061);
   ix3060 : mux21 port map ( Y=>nx3059, A0=>nx2963, A1=>nx2971, S0=>nx2967);
   ix3062 : xnor2 port map ( Y=>nx3061, A0=>nx3063, A1=>nx3065);
   ix3064 : nand02 port map ( Y=>nx3063, A0=>nx5476, A1=>nx362);
   ix3066 : xnor2 port map ( Y=>nx3065, A0=>nx3067, A1=>nx3069);
   ix3068 : mux21 port map ( Y=>nx3067, A0=>nx2973, A1=>nx2979, S0=>nx2975);
   ix3070 : xnor2 port map ( Y=>nx3069, A0=>nx3071, A1=>nx3073);
   ix3072 : nand02 port map ( Y=>nx3071, A0=>nx5472, A1=>nx338);
   ix3074 : xnor2 port map ( Y=>nx3073, A0=>nx3075, A1=>nx3077);
   ix3076 : mux21 port map ( Y=>nx3075, A0=>nx2981, A1=>nx2987, S0=>nx2983);
   ix3078 : xnor2 port map ( Y=>nx3077, A0=>nx3079, A1=>nx3081);
   ix3080 : nand02 port map ( Y=>nx3079, A0=>nx5468, A1=>nx314);
   ix3082 : xnor2 port map ( Y=>nx3081, A0=>nx3083, A1=>nx3085);
   ix3084 : mux21 port map ( Y=>nx3083, A0=>nx2989, A1=>nx2995, S0=>nx2991);
   ix3086 : xnor2 port map ( Y=>nx3085, A0=>nx3087, A1=>nx3089);
   ix3088 : nand02 port map ( Y=>nx3087, A0=>nx5456, A1=>nx290);
   ix3090 : nand02 port map ( Y=>nx3089, A0=>nx5448, A1=>nx266);
   ix267 : mux21 port map ( Y=>nx266, A0=>C(8), A1=>lfsr_C_8, S0=>test_mode
   );
   ix2021 : nor03 port map ( Y=>nx2020, A0=>nx3033, A1=>nx5536, A2=>nx3095);
   ix4371 : nor02ii port map ( Y=>mac_output(9), A0=>RST, A1=>nx4366);
   ix4367 : nor02 port map ( Y=>nx4366, A0=>RST, A1=>nx3103);
   ix3104 : xnor2 port map ( Y=>nx3103, A0=>nx3105, A1=>nx3111);
   ix3106 : xnor2 port map ( Y=>nx3105, A0=>mac_unit_tempP_9, A1=>nx3860);
   mac_unit_MR_reg_Q_9 : dffr port map ( Q=>mac_unit_tempP_9, QB=>OPEN, D=>
      nx3848, CLK=>CLK, R=>RST);
   ix3112 : aoi22 port map ( Y=>nx3111, A0=>nx3836, A1=>mac_unit_tempP_8, B0
      =>nx1923, B1=>nx3822);
   ix3861 : aoi21 port map ( Y=>nx3860, A0=>nx3121, A1=>nx3125, B0=>nx2242);
   ix2089 : mux21 port map ( Y=>nx2088, A0=>B(9), A1=>lfsr_C_6, S0=>
      test_mode);
   ix3126 : xnor2 port map ( Y=>nx3125, A0=>nx2020, A1=>nx2010);
   ix2011 : xnor2 port map ( Y=>nx2010, A0=>nx3129, A1=>nx2006);
   ix2007 : xnor2 port map ( Y=>nx2006, A0=>nx1802, A1=>nx3135);
   ix1803 : mux21 port map ( Y=>nx1802, A0=>nx1784, A1=>nx1798, S0=>nx1788);
   ix3136 : xnor2 port map ( Y=>nx3135, A0=>nx3137, A1=>nx3139);
   ix3138 : nand02 port map ( Y=>nx3137, A0=>nx410, A1=>nx5488);
   ix3140 : xnor2 port map ( Y=>nx3139, A0=>nx3141, A1=>nx3145);
   ix3142 : mux21 port map ( Y=>nx3141, A0=>nx3143, A1=>nx3047, S0=>nx3043);
   ix3146 : xnor2 port map ( Y=>nx3145, A0=>nx3147, A1=>nx3149);
   ix3148 : nand02 port map ( Y=>nx3147, A0=>nx386, A1=>nx5484);
   ix3150 : xnor2 port map ( Y=>nx3149, A0=>nx3151, A1=>nx3153);
   ix3152 : mux21 port map ( Y=>nx3151, A0=>nx3049, A1=>nx3057, S0=>nx3053);
   ix3154 : xnor2 port map ( Y=>nx3153, A0=>nx3155, A1=>nx3157);
   ix3156 : nand02 port map ( Y=>nx3155, A0=>nx362, A1=>nx5480);
   ix3158 : xnor2 port map ( Y=>nx3157, A0=>nx3159, A1=>nx3161);
   ix3160 : mux21 port map ( Y=>nx3159, A0=>nx3059, A1=>nx3065, S0=>nx3061);
   ix3162 : xnor2 port map ( Y=>nx3161, A0=>nx3163, A1=>nx3165);
   ix3164 : nand02 port map ( Y=>nx3163, A0=>nx5476, A1=>nx338);
   ix3166 : xnor2 port map ( Y=>nx3165, A0=>nx3167, A1=>nx3169);
   ix3168 : mux21 port map ( Y=>nx3167, A0=>nx3067, A1=>nx3073, S0=>nx3069);
   ix3170 : xnor2 port map ( Y=>nx3169, A0=>nx3171, A1=>nx3173);
   ix3172 : nand02 port map ( Y=>nx3171, A0=>nx5472, A1=>nx314);
   ix3174 : xnor2 port map ( Y=>nx3173, A0=>nx3175, A1=>nx3177);
   ix3176 : mux21 port map ( Y=>nx3175, A0=>nx3075, A1=>nx3081, S0=>nx3077);
   ix3178 : xnor2 port map ( Y=>nx3177, A0=>nx3179, A1=>nx3181);
   ix3180 : nand02 port map ( Y=>nx3179, A0=>nx5468, A1=>nx290);
   ix3182 : xnor2 port map ( Y=>nx3181, A0=>nx3183, A1=>nx3185);
   ix3184 : mux21 port map ( Y=>nx3183, A0=>nx3083, A1=>nx3089, S0=>nx3085);
   ix3186 : xnor2 port map ( Y=>nx3185, A0=>nx3187, A1=>nx3189);
   ix3188 : nand02 port map ( Y=>nx3187, A0=>nx5456, A1=>nx266);
   ix3190 : nand02 port map ( Y=>nx3189, A0=>nx5448, A1=>nx242);
   ix243 : mux21 port map ( Y=>nx242, A0=>C(9), A1=>lfsr_C_9, S0=>test_mode
   );
   ix2243 : nor03 port map ( Y=>nx2242, A0=>nx3125, A1=>nx5536, A2=>nx3195);
   ix4379 : nor02ii port map ( Y=>mac_output(10), A0=>RST, A1=>nx4374);
   ix4375 : nor02 port map ( Y=>nx4374, A0=>RST, A1=>nx3203);
   ix3204 : xnor2 port map ( Y=>nx3203, A0=>nx3205, A1=>nx3211);
   ix3206 : xnor2 port map ( Y=>nx3205, A0=>mac_unit_tempP_10, A1=>nx3884);
   mac_unit_MR_reg_Q_10 : dffr port map ( Q=>mac_unit_tempP_10, QB=>OPEN, D
      =>nx3872, CLK=>CLK, R=>RST);
   ix3212 : aoi22 port map ( Y=>nx3211, A0=>nx3860, A1=>mac_unit_tempP_9, B0
      =>nx1922, B1=>nx3846);
   ix3885 : aoi21 port map ( Y=>nx3884, A0=>nx3221, A1=>nx3225, B0=>nx2464);
   ix2311 : mux21 port map ( Y=>nx2310, A0=>B(10), A1=>lfsr_C_5, S0=>
      test_mode);
   ix3226 : xnor2 port map ( Y=>nx3225, A0=>nx2242, A1=>nx2232);
   ix2233 : xnor2 port map ( Y=>nx2232, A0=>nx3229, A1=>nx2228);
   ix2229 : xnor2 port map ( Y=>nx2228, A0=>nx2024, A1=>nx3235);
   ix2025 : mux21 port map ( Y=>nx2024, A0=>nx2006, A1=>nx2020, S0=>nx2010);
   ix3236 : xnor2 port map ( Y=>nx3235, A0=>nx3237, A1=>nx3239);
   ix3238 : nand02 port map ( Y=>nx3237, A0=>nx410, A1=>nx5492);
   ix3240 : xnor2 port map ( Y=>nx3239, A0=>nx3241, A1=>nx3245);
   ix3242 : mux21 port map ( Y=>nx3241, A0=>nx3243, A1=>nx3139, S0=>nx3135);
   ix3246 : xnor2 port map ( Y=>nx3245, A0=>nx3247, A1=>nx3249);
   ix3248 : nand02 port map ( Y=>nx3247, A0=>nx386, A1=>nx5488);
   ix3250 : xnor2 port map ( Y=>nx3249, A0=>nx3251, A1=>nx3253);
   ix3252 : mux21 port map ( Y=>nx3251, A0=>nx3141, A1=>nx3149, S0=>nx3145);
   ix3254 : xnor2 port map ( Y=>nx3253, A0=>nx3255, A1=>nx3257);
   ix3256 : nand02 port map ( Y=>nx3255, A0=>nx362, A1=>nx5484);
   ix3258 : xnor2 port map ( Y=>nx3257, A0=>nx3259, A1=>nx3261);
   ix3260 : mux21 port map ( Y=>nx3259, A0=>nx3151, A1=>nx3157, S0=>nx3153);
   ix3262 : xnor2 port map ( Y=>nx3261, A0=>nx3263, A1=>nx3265);
   ix3264 : nand02 port map ( Y=>nx3263, A0=>nx5480, A1=>nx338);
   ix3266 : xnor2 port map ( Y=>nx3265, A0=>nx3267, A1=>nx3269);
   ix3268 : mux21 port map ( Y=>nx3267, A0=>nx3159, A1=>nx3165, S0=>nx3161);
   ix3270 : xnor2 port map ( Y=>nx3269, A0=>nx3271, A1=>nx3273);
   ix3272 : nand02 port map ( Y=>nx3271, A0=>nx5476, A1=>nx314);
   ix3274 : xnor2 port map ( Y=>nx3273, A0=>nx3275, A1=>nx3277);
   ix3276 : mux21 port map ( Y=>nx3275, A0=>nx3167, A1=>nx3173, S0=>nx3169);
   ix3278 : xnor2 port map ( Y=>nx3277, A0=>nx3279, A1=>nx3281);
   ix3280 : nand02 port map ( Y=>nx3279, A0=>nx5472, A1=>nx290);
   ix3282 : xnor2 port map ( Y=>nx3281, A0=>nx3283, A1=>nx3285);
   ix3284 : mux21 port map ( Y=>nx3283, A0=>nx3175, A1=>nx3181, S0=>nx3177);
   ix3286 : xnor2 port map ( Y=>nx3285, A0=>nx3287, A1=>nx3289);
   ix3288 : nand02 port map ( Y=>nx3287, A0=>nx5468, A1=>nx266);
   ix3290 : xnor2 port map ( Y=>nx3289, A0=>nx3291, A1=>nx3293);
   ix3292 : mux21 port map ( Y=>nx3291, A0=>nx3183, A1=>nx3189, S0=>nx3185);
   ix3294 : xnor2 port map ( Y=>nx3293, A0=>nx3295, A1=>nx3297);
   ix3296 : nand02 port map ( Y=>nx3295, A0=>nx5456, A1=>nx242);
   ix3298 : nand02 port map ( Y=>nx3297, A0=>nx5448, A1=>nx218);
   ix219 : mux21 port map ( Y=>nx218, A0=>C(10), A1=>lfsr_C_10, S0=>
      test_mode);
   ix2465 : nor03 port map ( Y=>nx2464, A0=>nx3225, A1=>nx5536, A2=>nx3303);
   ix4387 : nor02ii port map ( Y=>mac_output(11), A0=>RST, A1=>nx4382);
   ix4383 : nor02 port map ( Y=>nx4382, A0=>RST, A1=>nx3311);
   ix3312 : xnor2 port map ( Y=>nx3311, A0=>nx3313, A1=>nx3319);
   ix3314 : xnor2 port map ( Y=>nx3313, A0=>mac_unit_tempP_11, A1=>nx3908);
   mac_unit_MR_reg_Q_11 : dffr port map ( Q=>mac_unit_tempP_11, QB=>OPEN, D
      =>nx3896, CLK=>CLK, R=>RST);
   ix3320 : aoi22 port map ( Y=>nx3319, A0=>nx3884, A1=>mac_unit_tempP_10, 
      B0=>nx1921, B1=>nx3870);
   ix3909 : aoi21 port map ( Y=>nx3908, A0=>nx3329, A1=>nx3333, B0=>nx2686);
   ix2533 : mux21 port map ( Y=>nx2532, A0=>B(11), A1=>lfsr_C_4, S0=>
      test_mode);
   ix3334 : xnor2 port map ( Y=>nx3333, A0=>nx2464, A1=>nx2454);
   ix2455 : xnor2 port map ( Y=>nx2454, A0=>nx3337, A1=>nx2450);
   ix2451 : xnor2 port map ( Y=>nx2450, A0=>nx2246, A1=>nx3343);
   ix2247 : mux21 port map ( Y=>nx2246, A0=>nx2228, A1=>nx2242, S0=>nx2232);
   ix3344 : xnor2 port map ( Y=>nx3343, A0=>nx3345, A1=>nx3347);
   ix3346 : nand02 port map ( Y=>nx3345, A0=>nx410, A1=>nx5496);
   ix3348 : xnor2 port map ( Y=>nx3347, A0=>nx3349, A1=>nx3353);
   ix3350 : mux21 port map ( Y=>nx3349, A0=>nx3351, A1=>nx3239, S0=>nx3235);
   ix3354 : xnor2 port map ( Y=>nx3353, A0=>nx3355, A1=>nx3357);
   ix3356 : nand02 port map ( Y=>nx3355, A0=>nx386, A1=>nx5492);
   ix3358 : xnor2 port map ( Y=>nx3357, A0=>nx3359, A1=>nx3361);
   ix3360 : mux21 port map ( Y=>nx3359, A0=>nx3241, A1=>nx3249, S0=>nx3245);
   ix3362 : xnor2 port map ( Y=>nx3361, A0=>nx3363, A1=>nx3365);
   ix3364 : nand02 port map ( Y=>nx3363, A0=>nx362, A1=>nx5488);
   ix3366 : xnor2 port map ( Y=>nx3365, A0=>nx3367, A1=>nx3369);
   ix3368 : mux21 port map ( Y=>nx3367, A0=>nx3251, A1=>nx3257, S0=>nx3253);
   ix3370 : xnor2 port map ( Y=>nx3369, A0=>nx3371, A1=>nx3373);
   ix3372 : nand02 port map ( Y=>nx3371, A0=>nx338, A1=>nx5484);
   ix3374 : xnor2 port map ( Y=>nx3373, A0=>nx3375, A1=>nx3377);
   ix3376 : mux21 port map ( Y=>nx3375, A0=>nx3259, A1=>nx3265, S0=>nx3261);
   ix3378 : xnor2 port map ( Y=>nx3377, A0=>nx3379, A1=>nx3381);
   ix3380 : nand02 port map ( Y=>nx3379, A0=>nx5480, A1=>nx314);
   ix3382 : xnor2 port map ( Y=>nx3381, A0=>nx3383, A1=>nx3385);
   ix3384 : mux21 port map ( Y=>nx3383, A0=>nx3267, A1=>nx3273, S0=>nx3269);
   ix3386 : xnor2 port map ( Y=>nx3385, A0=>nx3387, A1=>nx3389);
   ix3388 : nand02 port map ( Y=>nx3387, A0=>nx5476, A1=>nx290);
   ix3390 : xnor2 port map ( Y=>nx3389, A0=>nx3391, A1=>nx3393);
   ix3392 : mux21 port map ( Y=>nx3391, A0=>nx3275, A1=>nx3281, S0=>nx3277);
   ix3394 : xnor2 port map ( Y=>nx3393, A0=>nx3395, A1=>nx3397);
   ix3396 : nand02 port map ( Y=>nx3395, A0=>nx5472, A1=>nx266);
   ix3398 : xnor2 port map ( Y=>nx3397, A0=>nx3399, A1=>nx3401);
   ix3400 : mux21 port map ( Y=>nx3399, A0=>nx3283, A1=>nx3289, S0=>nx3285);
   ix3402 : xnor2 port map ( Y=>nx3401, A0=>nx3403, A1=>nx3405);
   ix3404 : nand02 port map ( Y=>nx3403, A0=>nx5468, A1=>nx242);
   ix3406 : xnor2 port map ( Y=>nx3405, A0=>nx3407, A1=>nx3409);
   ix3408 : mux21 port map ( Y=>nx3407, A0=>nx3291, A1=>nx3297, S0=>nx3293);
   ix3410 : xnor2 port map ( Y=>nx3409, A0=>nx3411, A1=>nx3413);
   ix3412 : nand02 port map ( Y=>nx3411, A0=>nx5456, A1=>nx218);
   ix3414 : nand02 port map ( Y=>nx3413, A0=>nx5448, A1=>nx194);
   ix195 : mux21 port map ( Y=>nx194, A0=>C(11), A1=>lfsr_C_11, S0=>
      test_mode);
   ix2687 : nor03 port map ( Y=>nx2686, A0=>nx3333, A1=>nx5536, A2=>nx3417);
   ix4395 : nor02ii port map ( Y=>mac_output(12), A0=>RST, A1=>nx4390);
   ix4391 : nor02 port map ( Y=>nx4390, A0=>RST, A1=>nx3425);
   ix3426 : xnor2 port map ( Y=>nx3425, A0=>nx3427, A1=>nx3433);
   ix3428 : xnor2 port map ( Y=>nx3427, A0=>mac_unit_tempP_12, A1=>nx3932);
   mac_unit_MR_reg_Q_12 : dffr port map ( Q=>mac_unit_tempP_12, QB=>OPEN, D
      =>nx3920, CLK=>CLK, R=>RST);
   ix3434 : aoi22 port map ( Y=>nx3433, A0=>nx3908, A1=>mac_unit_tempP_11, 
      B0=>nx1919, B1=>nx3894);
   ix3933 : aoi21 port map ( Y=>nx3932, A0=>nx3443, A1=>nx3447, B0=>nx2908);
   ix2755 : mux21 port map ( Y=>nx2754, A0=>B(12), A1=>lfsr_C_3, S0=>
      test_mode);
   ix3448 : xnor2 port map ( Y=>nx3447, A0=>nx2686, A1=>nx2676);
   ix2677 : xnor2 port map ( Y=>nx2676, A0=>nx3451, A1=>nx2672);
   ix2673 : xnor2 port map ( Y=>nx2672, A0=>nx2468, A1=>nx3457);
   ix2469 : mux21 port map ( Y=>nx2468, A0=>nx2450, A1=>nx2464, S0=>nx2454);
   ix3458 : xnor2 port map ( Y=>nx3457, A0=>nx3459, A1=>nx3461);
   ix3460 : nand02 port map ( Y=>nx3459, A0=>nx410, A1=>nx5500);
   ix3462 : xnor2 port map ( Y=>nx3461, A0=>nx3463, A1=>nx3467);
   ix3464 : mux21 port map ( Y=>nx3463, A0=>nx3465, A1=>nx3347, S0=>nx3343);
   ix3468 : xnor2 port map ( Y=>nx3467, A0=>nx3469, A1=>nx3471);
   ix3470 : nand02 port map ( Y=>nx3469, A0=>nx386, A1=>nx5496);
   ix3472 : xnor2 port map ( Y=>nx3471, A0=>nx3473, A1=>nx3475);
   ix3474 : mux21 port map ( Y=>nx3473, A0=>nx3349, A1=>nx3357, S0=>nx3353);
   ix3476 : xnor2 port map ( Y=>nx3475, A0=>nx3477, A1=>nx3479);
   ix3478 : nand02 port map ( Y=>nx3477, A0=>nx362, A1=>nx5492);
   ix3480 : xnor2 port map ( Y=>nx3479, A0=>nx3481, A1=>nx3483);
   ix3482 : mux21 port map ( Y=>nx3481, A0=>nx3359, A1=>nx3365, S0=>nx3361);
   ix3484 : xnor2 port map ( Y=>nx3483, A0=>nx3485, A1=>nx3487);
   ix3486 : nand02 port map ( Y=>nx3485, A0=>nx338, A1=>nx5488);
   ix3488 : xnor2 port map ( Y=>nx3487, A0=>nx3489, A1=>nx3491);
   ix3490 : mux21 port map ( Y=>nx3489, A0=>nx3367, A1=>nx3373, S0=>nx3369);
   ix3492 : xnor2 port map ( Y=>nx3491, A0=>nx3493, A1=>nx3495);
   ix3494 : nand02 port map ( Y=>nx3493, A0=>nx5484, A1=>nx314);
   ix3496 : xnor2 port map ( Y=>nx3495, A0=>nx3497, A1=>nx3499);
   ix3498 : mux21 port map ( Y=>nx3497, A0=>nx3375, A1=>nx3381, S0=>nx3377);
   ix3500 : xnor2 port map ( Y=>nx3499, A0=>nx3501, A1=>nx3503);
   ix3502 : nand02 port map ( Y=>nx3501, A0=>nx5480, A1=>nx290);
   ix3504 : xnor2 port map ( Y=>nx3503, A0=>nx3505, A1=>nx3507);
   ix3506 : mux21 port map ( Y=>nx3505, A0=>nx3383, A1=>nx3389, S0=>nx3385);
   ix3508 : xnor2 port map ( Y=>nx3507, A0=>nx3509, A1=>nx3511);
   ix3510 : nand02 port map ( Y=>nx3509, A0=>nx5476, A1=>nx266);
   ix3512 : xnor2 port map ( Y=>nx3511, A0=>nx3513, A1=>nx3515);
   ix3514 : mux21 port map ( Y=>nx3513, A0=>nx3391, A1=>nx3397, S0=>nx3393);
   ix3516 : xnor2 port map ( Y=>nx3515, A0=>nx3517, A1=>nx3519);
   ix3518 : nand02 port map ( Y=>nx3517, A0=>nx5472, A1=>nx242);
   ix3520 : xnor2 port map ( Y=>nx3519, A0=>nx3521, A1=>nx3523);
   ix3522 : mux21 port map ( Y=>nx3521, A0=>nx3399, A1=>nx3405, S0=>nx3401);
   ix3524 : xnor2 port map ( Y=>nx3523, A0=>nx3525, A1=>nx3527);
   ix3526 : nand02 port map ( Y=>nx3525, A0=>nx5468, A1=>nx218);
   ix3528 : xnor2 port map ( Y=>nx3527, A0=>nx3529, A1=>nx3531);
   ix3530 : mux21 port map ( Y=>nx3529, A0=>nx3407, A1=>nx3413, S0=>nx3409);
   ix3532 : xnor2 port map ( Y=>nx3531, A0=>nx3533, A1=>nx3535);
   ix3534 : nand02 port map ( Y=>nx3533, A0=>nx5456, A1=>nx194);
   ix3536 : nand02 port map ( Y=>nx3535, A0=>nx5448, A1=>nx170);
   ix171 : mux21 port map ( Y=>nx170, A0=>C(12), A1=>lfsr_C_12, S0=>
      test_mode);
   ix2909 : nor03 port map ( Y=>nx2908, A0=>nx3447, A1=>nx5536, A2=>nx3541);
   ix4403 : nor02ii port map ( Y=>mac_output(13), A0=>RST, A1=>nx4398);
   ix4399 : nor02 port map ( Y=>nx4398, A0=>RST, A1=>nx3549);
   ix3550 : xnor2 port map ( Y=>nx3549, A0=>nx3551, A1=>nx3557);
   ix3552 : xnor2 port map ( Y=>nx3551, A0=>mac_unit_tempP_13, A1=>nx3956);
   mac_unit_MR_reg_Q_13 : dffr port map ( Q=>mac_unit_tempP_13, QB=>OPEN, D
      =>nx3944, CLK=>CLK, R=>RST);
   ix3558 : aoi22 port map ( Y=>nx3557, A0=>nx3932, A1=>mac_unit_tempP_12, 
      B0=>nx1917, B1=>nx3918);
   ix3957 : aoi21 port map ( Y=>nx3956, A0=>nx3567, A1=>nx3571, B0=>nx3130);
   ix2977 : mux21 port map ( Y=>nx2976, A0=>B(13), A1=>lfsr_C_2, S0=>
      test_mode);
   ix3572 : xnor2 port map ( Y=>nx3571, A0=>nx2908, A1=>nx2898);
   ix2899 : xnor2 port map ( Y=>nx2898, A0=>nx3575, A1=>nx2894);
   ix2895 : xnor2 port map ( Y=>nx2894, A0=>nx2690, A1=>nx3581);
   ix2691 : mux21 port map ( Y=>nx2690, A0=>nx2672, A1=>nx2686, S0=>nx2676);
   ix3582 : xnor2 port map ( Y=>nx3581, A0=>nx3583, A1=>nx3585);
   ix3584 : nand02 port map ( Y=>nx3583, A0=>nx410, A1=>nx5504);
   ix3586 : xnor2 port map ( Y=>nx3585, A0=>nx3587, A1=>nx3591);
   ix3588 : mux21 port map ( Y=>nx3587, A0=>nx3589, A1=>nx3461, S0=>nx3457);
   ix3592 : xnor2 port map ( Y=>nx3591, A0=>nx3593, A1=>nx3595);
   ix3594 : nand02 port map ( Y=>nx3593, A0=>nx386, A1=>nx5500);
   ix3596 : xnor2 port map ( Y=>nx3595, A0=>nx3597, A1=>nx3599);
   ix3598 : mux21 port map ( Y=>nx3597, A0=>nx3463, A1=>nx3471, S0=>nx3467);
   ix3600 : xnor2 port map ( Y=>nx3599, A0=>nx3601, A1=>nx3603);
   ix3602 : nand02 port map ( Y=>nx3601, A0=>nx362, A1=>nx5496);
   ix3604 : xnor2 port map ( Y=>nx3603, A0=>nx3605, A1=>nx3607);
   ix3606 : mux21 port map ( Y=>nx3605, A0=>nx3473, A1=>nx3479, S0=>nx3475);
   ix3608 : xnor2 port map ( Y=>nx3607, A0=>nx3609, A1=>nx3611);
   ix3610 : nand02 port map ( Y=>nx3609, A0=>nx338, A1=>nx5492);
   ix3612 : xnor2 port map ( Y=>nx3611, A0=>nx3613, A1=>nx3615);
   ix3614 : mux21 port map ( Y=>nx3613, A0=>nx3481, A1=>nx3487, S0=>nx3483);
   ix3616 : xnor2 port map ( Y=>nx3615, A0=>nx3617, A1=>nx3619);
   ix3618 : nand02 port map ( Y=>nx3617, A0=>nx314, A1=>nx5488);
   ix3620 : xnor2 port map ( Y=>nx3619, A0=>nx3621, A1=>nx3623);
   ix3622 : mux21 port map ( Y=>nx3621, A0=>nx3489, A1=>nx3495, S0=>nx3491);
   ix3624 : xnor2 port map ( Y=>nx3623, A0=>nx3625, A1=>nx3627);
   ix3626 : nand02 port map ( Y=>nx3625, A0=>nx5484, A1=>nx290);
   ix3628 : xnor2 port map ( Y=>nx3627, A0=>nx3629, A1=>nx3631);
   ix3630 : mux21 port map ( Y=>nx3629, A0=>nx3497, A1=>nx3503, S0=>nx3499);
   ix3632 : xnor2 port map ( Y=>nx3631, A0=>nx3633, A1=>nx3635);
   ix3634 : nand02 port map ( Y=>nx3633, A0=>nx5480, A1=>nx266);
   ix3636 : xnor2 port map ( Y=>nx3635, A0=>nx3637, A1=>nx3639);
   ix3638 : mux21 port map ( Y=>nx3637, A0=>nx3505, A1=>nx3511, S0=>nx3507);
   ix3640 : xnor2 port map ( Y=>nx3639, A0=>nx3641, A1=>nx3643);
   ix3642 : nand02 port map ( Y=>nx3641, A0=>nx5476, A1=>nx242);
   ix3644 : xnor2 port map ( Y=>nx3643, A0=>nx3645, A1=>nx3647);
   ix3646 : mux21 port map ( Y=>nx3645, A0=>nx3513, A1=>nx3519, S0=>nx3515);
   ix3648 : xnor2 port map ( Y=>nx3647, A0=>nx3649, A1=>nx3651);
   ix3650 : nand02 port map ( Y=>nx3649, A0=>nx5472, A1=>nx218);
   ix3652 : xnor2 port map ( Y=>nx3651, A0=>nx3653, A1=>nx3655);
   ix3654 : mux21 port map ( Y=>nx3653, A0=>nx3521, A1=>nx3527, S0=>nx3523);
   ix3656 : xnor2 port map ( Y=>nx3655, A0=>nx3657, A1=>nx3659);
   ix3658 : nand02 port map ( Y=>nx3657, A0=>nx5468, A1=>nx194);
   ix3660 : xnor2 port map ( Y=>nx3659, A0=>nx3661, A1=>nx3663);
   ix3662 : mux21 port map ( Y=>nx3661, A0=>nx3529, A1=>nx3535, S0=>nx3531);
   ix3664 : xnor2 port map ( Y=>nx3663, A0=>nx3665, A1=>nx3667);
   ix3666 : nand02 port map ( Y=>nx3665, A0=>nx5456, A1=>nx170);
   ix3668 : nand02 port map ( Y=>nx3667, A0=>nx5448, A1=>nx146);
   ix147 : mux21 port map ( Y=>nx146, A0=>C(13), A1=>lfsr_C_13, S0=>
      test_mode);
   ix3131 : nor03 port map ( Y=>nx3130, A0=>nx3571, A1=>nx5536, A2=>nx3673);
   ix4411 : nor02ii port map ( Y=>mac_output(14), A0=>RST, A1=>nx4406);
   ix4407 : nor02 port map ( Y=>nx4406, A0=>RST, A1=>nx3681);
   ix3682 : xnor2 port map ( Y=>nx3681, A0=>nx3683, A1=>nx3687);
   ix3684 : xnor2 port map ( Y=>nx3683, A0=>mac_unit_tempP_14, A1=>nx3980);
   mac_unit_MR_reg_Q_14 : dffr port map ( Q=>mac_unit_tempP_14, QB=>OPEN, D
      =>nx3968, CLK=>CLK, R=>RST);
   ix3688 : aoi22 port map ( Y=>nx3687, A0=>nx3956, A1=>mac_unit_tempP_13, 
      B0=>nx1915, B1=>nx3942);
   ix3981 : aoi21 port map ( Y=>nx3980, A0=>nx3697, A1=>nx3701, B0=>nx3352);
   ix3199 : mux21 port map ( Y=>nx3198, A0=>B(14), A1=>lfsr_C_1, S0=>
      test_mode);
   ix3702 : xnor2 port map ( Y=>nx3701, A0=>nx3130, A1=>nx3120);
   ix3121 : xnor2 port map ( Y=>nx3120, A0=>nx3705, A1=>nx3116);
   ix3117 : xnor2 port map ( Y=>nx3116, A0=>nx2912, A1=>nx3709);
   ix2913 : mux21 port map ( Y=>nx2912, A0=>nx2894, A1=>nx2908, S0=>nx2898);
   ix3710 : xnor2 port map ( Y=>nx3709, A0=>nx3711, A1=>nx3713);
   ix3712 : nand02 port map ( Y=>nx3711, A0=>nx410, A1=>nx5508);
   ix3714 : xnor2 port map ( Y=>nx3713, A0=>nx3715, A1=>nx3719);
   ix3716 : mux21 port map ( Y=>nx3715, A0=>nx3717, A1=>nx3585, S0=>nx3581);
   ix3720 : xnor2 port map ( Y=>nx3719, A0=>nx3721, A1=>nx3723);
   ix3722 : nand02 port map ( Y=>nx3721, A0=>nx386, A1=>nx5504);
   ix3724 : xnor2 port map ( Y=>nx3723, A0=>nx3725, A1=>nx3727);
   ix3726 : mux21 port map ( Y=>nx3725, A0=>nx3587, A1=>nx3595, S0=>nx3591);
   ix3728 : xnor2 port map ( Y=>nx3727, A0=>nx3729, A1=>nx3731);
   ix3730 : nand02 port map ( Y=>nx3729, A0=>nx362, A1=>nx5500);
   ix3732 : xnor2 port map ( Y=>nx3731, A0=>nx3733, A1=>nx3735);
   ix3734 : mux21 port map ( Y=>nx3733, A0=>nx3597, A1=>nx3603, S0=>nx3599);
   ix3736 : xnor2 port map ( Y=>nx3735, A0=>nx3737, A1=>nx3739);
   ix3738 : nand02 port map ( Y=>nx3737, A0=>nx338, A1=>nx5496);
   ix3740 : xnor2 port map ( Y=>nx3739, A0=>nx3741, A1=>nx3743);
   ix3742 : mux21 port map ( Y=>nx3741, A0=>nx3605, A1=>nx3611, S0=>nx3607);
   ix3744 : xnor2 port map ( Y=>nx3743, A0=>nx3745, A1=>nx3747);
   ix3746 : nand02 port map ( Y=>nx3745, A0=>nx314, A1=>nx5492);
   ix3748 : xnor2 port map ( Y=>nx3747, A0=>nx3749, A1=>nx3751);
   ix3750 : mux21 port map ( Y=>nx3749, A0=>nx3613, A1=>nx3619, S0=>nx3615);
   ix3752 : xnor2 port map ( Y=>nx3751, A0=>nx3753, A1=>nx3755);
   ix3754 : nand02 port map ( Y=>nx3753, A0=>nx5488, A1=>nx290);
   ix3756 : xnor2 port map ( Y=>nx3755, A0=>nx3757, A1=>nx3759);
   ix3758 : mux21 port map ( Y=>nx3757, A0=>nx3621, A1=>nx3627, S0=>nx3623);
   ix3760 : xnor2 port map ( Y=>nx3759, A0=>nx3761, A1=>nx3763);
   ix3762 : nand02 port map ( Y=>nx3761, A0=>nx5484, A1=>nx266);
   ix3764 : xnor2 port map ( Y=>nx3763, A0=>nx3765, A1=>nx3767);
   ix3766 : mux21 port map ( Y=>nx3765, A0=>nx3629, A1=>nx3635, S0=>nx3631);
   ix3768 : xnor2 port map ( Y=>nx3767, A0=>nx3769, A1=>nx3771);
   ix3770 : nand02 port map ( Y=>nx3769, A0=>nx5480, A1=>nx242);
   ix3772 : xnor2 port map ( Y=>nx3771, A0=>nx3773, A1=>nx3775);
   ix3774 : mux21 port map ( Y=>nx3773, A0=>nx3637, A1=>nx3643, S0=>nx3639);
   ix3776 : xnor2 port map ( Y=>nx3775, A0=>nx3777, A1=>nx3779);
   ix3778 : nand02 port map ( Y=>nx3777, A0=>nx5476, A1=>nx218);
   ix3780 : xnor2 port map ( Y=>nx3779, A0=>nx3781, A1=>nx3783);
   ix3782 : mux21 port map ( Y=>nx3781, A0=>nx3645, A1=>nx3651, S0=>nx3647);
   ix3784 : xnor2 port map ( Y=>nx3783, A0=>nx3785, A1=>nx3787);
   ix3786 : nand02 port map ( Y=>nx3785, A0=>nx5472, A1=>nx194);
   ix3788 : xnor2 port map ( Y=>nx3787, A0=>nx3789, A1=>nx3791);
   ix3790 : mux21 port map ( Y=>nx3789, A0=>nx3653, A1=>nx3659, S0=>nx3655);
   ix3792 : xnor2 port map ( Y=>nx3791, A0=>nx3793, A1=>nx3795);
   ix3794 : nand02 port map ( Y=>nx3793, A0=>nx5468, A1=>nx170);
   ix3796 : xnor2 port map ( Y=>nx3795, A0=>nx3797, A1=>nx3799);
   ix3798 : mux21 port map ( Y=>nx3797, A0=>nx3661, A1=>nx3667, S0=>nx3663);
   ix3800 : xnor2 port map ( Y=>nx3799, A0=>nx3801, A1=>nx3803);
   ix3802 : nand02 port map ( Y=>nx3801, A0=>nx5456, A1=>nx146);
   ix3804 : nand02 port map ( Y=>nx3803, A0=>nx5450, A1=>nx122);
   ix123 : mux21 port map ( Y=>nx122, A0=>C(14), A1=>lfsr_C_14, S0=>
      test_mode);
   ix3353 : nor03 port map ( Y=>nx3352, A0=>nx3701, A1=>nx5536, A2=>nx3807);
   ix4419 : nor02ii port map ( Y=>mac_output(15), A0=>RST, A1=>nx4414);
   ix4415 : nor02 port map ( Y=>nx4414, A0=>RST, A1=>nx3815);
   ix3816 : xnor2 port map ( Y=>nx3815, A0=>nx3817, A1=>nx3823);
   ix3818 : xnor2 port map ( Y=>nx3817, A0=>mac_unit_tempP_15, A1=>nx4004);
   mac_unit_MR_reg_Q_15 : dffr port map ( Q=>mac_unit_tempP_15, QB=>OPEN, D
      =>nx3992, CLK=>CLK, R=>RST);
   ix3824 : aoi22 port map ( Y=>nx3823, A0=>nx3980, A1=>mac_unit_tempP_14, 
      B0=>nx1913, B1=>nx3966);
   ix4005 : aoi21 port map ( Y=>nx4004, A0=>nx3833, A1=>nx3837, B0=>nx3574);
   ix3421 : mux21 port map ( Y=>nx3420, A0=>B(15), A1=>lfsr_B_15, S0=>
      test_mode);
   ix3838 : xnor2 port map ( Y=>nx3837, A0=>nx3352, A1=>nx3342);
   ix3343 : xnor2 port map ( Y=>nx3342, A0=>nx3841, A1=>nx3338);
   ix3339 : xnor2 port map ( Y=>nx3338, A0=>nx3134, A1=>nx3847);
   ix3135 : mux21 port map ( Y=>nx3134, A0=>nx3116, A1=>nx3130, S0=>nx3120);
   ix3848 : xnor2 port map ( Y=>nx3847, A0=>nx3849, A1=>nx3851);
   ix3850 : nand02 port map ( Y=>nx3849, A0=>nx410, A1=>nx5512);
   ix3852 : xnor2 port map ( Y=>nx3851, A0=>nx3853, A1=>nx3857);
   ix3854 : mux21 port map ( Y=>nx3853, A0=>nx3855, A1=>nx3713, S0=>nx3709);
   ix3858 : xnor2 port map ( Y=>nx3857, A0=>nx3859, A1=>nx3861);
   ix3860 : nand02 port map ( Y=>nx3859, A0=>nx386, A1=>nx5508);
   ix3862 : xnor2 port map ( Y=>nx3861, A0=>nx3863, A1=>nx3865);
   ix3864 : mux21 port map ( Y=>nx3863, A0=>nx3715, A1=>nx3723, S0=>nx3719);
   ix3866 : xnor2 port map ( Y=>nx3865, A0=>nx3867, A1=>nx3869);
   ix3868 : nand02 port map ( Y=>nx3867, A0=>nx362, A1=>nx5504);
   ix3870 : xnor2 port map ( Y=>nx3869, A0=>nx3871, A1=>nx3873);
   ix3872 : mux21 port map ( Y=>nx3871, A0=>nx3725, A1=>nx3731, S0=>nx3727);
   ix3874 : xnor2 port map ( Y=>nx3873, A0=>nx3875, A1=>nx3877);
   ix3876 : nand02 port map ( Y=>nx3875, A0=>nx338, A1=>nx5500);
   ix3878 : xnor2 port map ( Y=>nx3877, A0=>nx3879, A1=>nx3881);
   ix3880 : mux21 port map ( Y=>nx3879, A0=>nx3733, A1=>nx3739, S0=>nx3735);
   ix3882 : xnor2 port map ( Y=>nx3881, A0=>nx3883, A1=>nx3885);
   ix3884 : nand02 port map ( Y=>nx3883, A0=>nx314, A1=>nx5496);
   ix3886 : xnor2 port map ( Y=>nx3885, A0=>nx3887, A1=>nx3889);
   ix3888 : mux21 port map ( Y=>nx3887, A0=>nx3741, A1=>nx3747, S0=>nx3743);
   ix3890 : xnor2 port map ( Y=>nx3889, A0=>nx3891, A1=>nx3893);
   ix3892 : nand02 port map ( Y=>nx3891, A0=>nx290, A1=>nx5492);
   ix3894 : xnor2 port map ( Y=>nx3893, A0=>nx3895, A1=>nx3897);
   ix3896 : mux21 port map ( Y=>nx3895, A0=>nx3749, A1=>nx3755, S0=>nx3751);
   ix3898 : xnor2 port map ( Y=>nx3897, A0=>nx3899, A1=>nx3901);
   ix3900 : nand02 port map ( Y=>nx3899, A0=>nx5488, A1=>nx266);
   ix3902 : xnor2 port map ( Y=>nx3901, A0=>nx3903, A1=>nx3905);
   ix3904 : mux21 port map ( Y=>nx3903, A0=>nx3757, A1=>nx3763, S0=>nx3759);
   ix3906 : xnor2 port map ( Y=>nx3905, A0=>nx3907, A1=>nx3909);
   ix3908 : nand02 port map ( Y=>nx3907, A0=>nx5484, A1=>nx242);
   ix3910 : xnor2 port map ( Y=>nx3909, A0=>nx3911, A1=>nx3913);
   ix3912 : mux21 port map ( Y=>nx3911, A0=>nx3765, A1=>nx3771, S0=>nx3767);
   ix3914 : xnor2 port map ( Y=>nx3913, A0=>nx3915, A1=>nx3917);
   ix3916 : nand02 port map ( Y=>nx3915, A0=>nx5480, A1=>nx218);
   ix3918 : xnor2 port map ( Y=>nx3917, A0=>nx3919, A1=>nx3921);
   ix3920 : mux21 port map ( Y=>nx3919, A0=>nx3773, A1=>nx3779, S0=>nx3775);
   ix3922 : xnor2 port map ( Y=>nx3921, A0=>nx3923, A1=>nx3925);
   ix3924 : nand02 port map ( Y=>nx3923, A0=>nx5476, A1=>nx194);
   ix3926 : xnor2 port map ( Y=>nx3925, A0=>nx3927, A1=>nx3929);
   ix3928 : mux21 port map ( Y=>nx3927, A0=>nx3781, A1=>nx3787, S0=>nx3783);
   ix3930 : xnor2 port map ( Y=>nx3929, A0=>nx3931, A1=>nx3933);
   ix3932 : nand02 port map ( Y=>nx3931, A0=>nx5472, A1=>nx170);
   ix3934 : xnor2 port map ( Y=>nx3933, A0=>nx3935, A1=>nx3937);
   ix3936 : mux21 port map ( Y=>nx3935, A0=>nx3789, A1=>nx3795, S0=>nx3791);
   ix3938 : xnor2 port map ( Y=>nx3937, A0=>nx3939, A1=>nx3941);
   ix3940 : nand02 port map ( Y=>nx3939, A0=>nx5468, A1=>nx146);
   ix3942 : xnor2 port map ( Y=>nx3941, A0=>nx3943, A1=>nx3945);
   ix3944 : mux21 port map ( Y=>nx3943, A0=>nx3797, A1=>nx3803, S0=>nx3799);
   ix3946 : xnor2 port map ( Y=>nx3945, A0=>nx3947, A1=>nx3949);
   ix3948 : nand02 port map ( Y=>nx3947, A0=>nx5456, A1=>nx122);
   ix99 : mux21 port map ( Y=>nx98, A0=>C(15), A1=>lfsr_C_15, S0=>test_mode
   );
   ix3575 : nor03 port map ( Y=>nx3574, A0=>nx3837, A1=>nx5536, A2=>nx3955);
   ix4427 : nor02ii port map ( Y=>mac_output(16), A0=>RST, A1=>nx4422);
   ix4423 : nor02 port map ( Y=>nx4422, A0=>RST, A1=>nx3963);
   ix3964 : xnor2 port map ( Y=>nx3963, A0=>nx3965, A1=>nx3971);
   ix3966 : xnor2 port map ( Y=>nx3965, A0=>mac_unit_tempP_16, A1=>nx4022);
   mac_unit_MR_reg_Q_16 : dffr port map ( Q=>mac_unit_tempP_16, QB=>OPEN, D
      =>nx4016, CLK=>CLK, R=>RST);
   ix3972 : aoi22 port map ( Y=>nx3971, A0=>nx4004, A1=>mac_unit_tempP_15, 
      B0=>nx1912, B1=>nx3990);
   ix4023 : xnor2 port map ( Y=>nx4022, A0=>nx3574, A1=>nx3979);
   ix3980 : xnor2 port map ( Y=>nx3979, A0=>nx3981, A1=>nx3983);
   ix3984 : xnor2 port map ( Y=>nx3983, A0=>nx3356, A1=>nx3332);
   ix3357 : mux21 port map ( Y=>nx3356, A0=>nx3338, A1=>nx3352, S0=>nx3342);
   ix3333 : xnor2 port map ( Y=>nx3332, A0=>nx3989, A1=>nx3328);
   ix3990 : nand02 port map ( Y=>nx3989, A0=>nx410, A1=>nx5516);
   ix3329 : xnor2 port map ( Y=>nx3328, A0=>nx3993, A1=>nx3100);
   ix3994 : mux21 port map ( Y=>nx3993, A0=>nx3995, A1=>nx3851, S0=>nx3847);
   ix3101 : xnor2 port map ( Y=>nx3100, A0=>nx3999, A1=>nx3096);
   ix4000 : nand02 port map ( Y=>nx3999, A0=>nx386, A1=>nx5512);
   ix3097 : xnor2 port map ( Y=>nx3096, A0=>nx4003, A1=>nx2868);
   ix4004 : mux21 port map ( Y=>nx4003, A0=>nx3853, A1=>nx3861, S0=>nx3857);
   ix2869 : xnor2 port map ( Y=>nx2868, A0=>nx4007, A1=>nx2864);
   ix4008 : nand02 port map ( Y=>nx4007, A0=>nx362, A1=>nx5508);
   ix2865 : xnor2 port map ( Y=>nx2864, A0=>nx4011, A1=>nx2636);
   ix4012 : mux21 port map ( Y=>nx4011, A0=>nx3863, A1=>nx3869, S0=>nx3865);
   ix2637 : xnor2 port map ( Y=>nx2636, A0=>nx4015, A1=>nx2632);
   ix4016 : nand02 port map ( Y=>nx4015, A0=>nx338, A1=>nx5504);
   ix2633 : xnor2 port map ( Y=>nx2632, A0=>nx4019, A1=>nx2404);
   ix4020 : mux21 port map ( Y=>nx4019, A0=>nx3871, A1=>nx3877, S0=>nx3873);
   ix2405 : xnor2 port map ( Y=>nx2404, A0=>nx4023, A1=>nx2400);
   ix4024 : nand02 port map ( Y=>nx4023, A0=>nx314, A1=>nx5500);
   ix2401 : xnor2 port map ( Y=>nx2400, A0=>nx4027, A1=>nx2172);
   ix4028 : mux21 port map ( Y=>nx4027, A0=>nx3879, A1=>nx3885, S0=>nx3881);
   ix2173 : xnor2 port map ( Y=>nx2172, A0=>nx4031, A1=>nx2168);
   ix4032 : nand02 port map ( Y=>nx4031, A0=>nx290, A1=>nx5496);
   ix2169 : xnor2 port map ( Y=>nx2168, A0=>nx4035, A1=>nx1940);
   ix4036 : mux21 port map ( Y=>nx4035, A0=>nx3887, A1=>nx3893, S0=>nx3889);
   ix1941 : xnor2 port map ( Y=>nx1940, A0=>nx4038, A1=>nx1936);
   ix4039 : nand02 port map ( Y=>nx4038, A0=>nx5492, A1=>nx266);
   ix1937 : xnor2 port map ( Y=>nx1936, A0=>nx4041, A1=>nx1708);
   ix4042 : mux21 port map ( Y=>nx4041, A0=>nx3895, A1=>nx3901, S0=>nx3897);
   ix1709 : xnor2 port map ( Y=>nx1708, A0=>nx4045, A1=>nx1704);
   ix4046 : nand02 port map ( Y=>nx4045, A0=>nx5488, A1=>nx242);
   ix1705 : xnor2 port map ( Y=>nx1704, A0=>nx4049, A1=>nx1476);
   ix4050 : mux21 port map ( Y=>nx4049, A0=>nx3903, A1=>nx3909, S0=>nx3905);
   ix1477 : xnor2 port map ( Y=>nx1476, A0=>nx4053, A1=>nx1472);
   ix4054 : nand02 port map ( Y=>nx4053, A0=>nx5484, A1=>nx218);
   ix1473 : xnor2 port map ( Y=>nx1472, A0=>nx4056, A1=>nx1244);
   ix4057 : mux21 port map ( Y=>nx4056, A0=>nx3911, A1=>nx3917, S0=>nx3913);
   ix1245 : xnor2 port map ( Y=>nx1244, A0=>nx4059, A1=>nx1240);
   ix4060 : nand02 port map ( Y=>nx4059, A0=>nx5480, A1=>nx194);
   ix1241 : xnor2 port map ( Y=>nx1240, A0=>nx4063, A1=>nx1012);
   ix4064 : mux21 port map ( Y=>nx4063, A0=>nx3919, A1=>nx3925, S0=>nx3921);
   ix1013 : xnor2 port map ( Y=>nx1012, A0=>nx4067, A1=>nx1008);
   ix4068 : nand02 port map ( Y=>nx4067, A0=>nx5476, A1=>nx170);
   ix1009 : xnor2 port map ( Y=>nx1008, A0=>nx4071, A1=>nx780);
   ix4072 : mux21 port map ( Y=>nx4071, A0=>nx3927, A1=>nx3933, S0=>nx3929);
   ix781 : xnor2 port map ( Y=>nx780, A0=>nx4074, A1=>nx776);
   ix4075 : nand02 port map ( Y=>nx4074, A0=>nx5472, A1=>nx146);
   ix777 : xnor2 port map ( Y=>nx776, A0=>nx4077, A1=>nx548);
   ix4078 : mux21 port map ( Y=>nx4077, A0=>nx3935, A1=>nx3941, S0=>nx3937);
   ix549 : xnor2 port map ( Y=>nx548, A0=>nx4081, A1=>nx544);
   ix4082 : nand02 port map ( Y=>nx4081, A0=>nx5468, A1=>nx122);
   ix545 : aoi21 port map ( Y=>nx544, A0=>nx4085, A1=>nx4087, B0=>nx520);
   ix4088 : mux21 port map ( Y=>nx4087, A0=>nx3943, A1=>nx3949, S0=>nx3945);
   ix521 : nor03 port map ( Y=>nx520, A0=>nx4087, A1=>nx2583, A2=>nx5550);
   ix4435 : nor02 port map ( Y=>mac_output(17), A0=>RST, A1=>nx4095);
   ix4096 : nand02 port map ( Y=>nx4095, A0=>nx2523, A1=>nx4034);
   ix4035 : xnor2 port map ( Y=>nx4034, A0=>nx1909, A1=>nx4239);
   ix4043 : xnor2 port map ( Y=>nx1909, A0=>mac_unit_tempP_17, A1=>nx4105);
   mac_unit_MR_reg_Q_17 : dffr port map ( Q=>mac_unit_tempP_17, QB=>OPEN, D
      =>nx4034, CLK=>CLK, R=>RST);
   ix4106 : xnor2 port map ( Y=>nx4105, A0=>nx4107, A1=>nx4111);
   ix4108 : mux21 port map ( Y=>nx4107, A0=>nx4109, A1=>nx3983, S0=>nx3979);
   ix4112 : xnor2 port map ( Y=>nx4111, A0=>nx4113, A1=>nx4115);
   ix4114 : nand02 port map ( Y=>nx4113, A0=>nx410, A1=>nx5520);
   ix4116 : xnor2 port map ( Y=>nx4115, A0=>nx3360, A1=>nx3322);
   ix3361 : mux21 port map ( Y=>nx3360, A0=>nx3328, A1=>nx3356, S0=>nx3332);
   ix3323 : xnor2 port map ( Y=>nx3322, A0=>nx4121, A1=>nx3318);
   ix4122 : nand02 port map ( Y=>nx4121, A0=>nx386, A1=>nx5516);
   ix3319 : xnor2 port map ( Y=>nx3318, A0=>nx4125, A1=>nx3090);
   ix4126 : mux21 port map ( Y=>nx4125, A0=>nx4127, A1=>nx3993, S0=>nx3100);
   ix3091 : xnor2 port map ( Y=>nx3090, A0=>nx4131, A1=>nx3086);
   ix4132 : nand02 port map ( Y=>nx4131, A0=>nx362, A1=>nx5512);
   ix3087 : xnor2 port map ( Y=>nx3086, A0=>nx4135, A1=>nx2858);
   ix4136 : mux21 port map ( Y=>nx4135, A0=>nx4137, A1=>nx4003, S0=>nx2868);
   ix2859 : xnor2 port map ( Y=>nx2858, A0=>nx4141, A1=>nx2854);
   ix4142 : nand02 port map ( Y=>nx4141, A0=>nx338, A1=>nx5508);
   ix2855 : xnor2 port map ( Y=>nx2854, A0=>nx4145, A1=>nx2626);
   ix4146 : mux21 port map ( Y=>nx4145, A0=>nx4147, A1=>nx4011, S0=>nx2636);
   ix2627 : xnor2 port map ( Y=>nx2626, A0=>nx4151, A1=>nx2622);
   ix4152 : nand02 port map ( Y=>nx4151, A0=>nx314, A1=>nx5504);
   ix2623 : xnor2 port map ( Y=>nx2622, A0=>nx4155, A1=>nx2394);
   ix4156 : mux21 port map ( Y=>nx4155, A0=>nx4157, A1=>nx4019, S0=>nx2404);
   ix2395 : xnor2 port map ( Y=>nx2394, A0=>nx4161, A1=>nx2390);
   ix4162 : nand02 port map ( Y=>nx4161, A0=>nx290, A1=>nx5500);
   ix2391 : xnor2 port map ( Y=>nx2390, A0=>nx4164, A1=>nx2162);
   ix4165 : mux21 port map ( Y=>nx4164, A0=>nx4167, A1=>nx4027, S0=>nx2172);
   ix2163 : xnor2 port map ( Y=>nx2162, A0=>nx4171, A1=>nx2158);
   ix4172 : nand02 port map ( Y=>nx4171, A0=>nx266, A1=>nx5496);
   ix2159 : xnor2 port map ( Y=>nx2158, A0=>nx4175, A1=>nx1930);
   ix4176 : mux21 port map ( Y=>nx4175, A0=>nx4177, A1=>nx4035, S0=>nx1940);
   ix1931 : xnor2 port map ( Y=>nx1930, A0=>nx4181, A1=>nx1926);
   ix4182 : nand02 port map ( Y=>nx4181, A0=>nx5492, A1=>nx242);
   ix1927 : xnor2 port map ( Y=>nx1926, A0=>nx4185, A1=>nx1698);
   ix4186 : mux21 port map ( Y=>nx4185, A0=>nx4187, A1=>nx4041, S0=>nx1708);
   ix1699 : xnor2 port map ( Y=>nx1698, A0=>nx4191, A1=>nx1694);
   ix4192 : nand02 port map ( Y=>nx4191, A0=>nx5488, A1=>nx218);
   ix1695 : xnor2 port map ( Y=>nx1694, A0=>nx4195, A1=>nx1466);
   ix4196 : mux21 port map ( Y=>nx4195, A0=>nx4197, A1=>nx4049, S0=>nx1476);
   ix1467 : xnor2 port map ( Y=>nx1466, A0=>nx4200, A1=>nx1462);
   ix4201 : nand02 port map ( Y=>nx4200, A0=>nx5484, A1=>nx194);
   ix1463 : xnor2 port map ( Y=>nx1462, A0=>nx4203, A1=>nx1234);
   ix4204 : mux21 port map ( Y=>nx4203, A0=>nx4205, A1=>nx4056, S0=>nx1244);
   ix1235 : xnor2 port map ( Y=>nx1234, A0=>nx4209, A1=>nx1230);
   ix4210 : nand02 port map ( Y=>nx4209, A0=>nx5480, A1=>nx170);
   ix1231 : xnor2 port map ( Y=>nx1230, A0=>nx4213, A1=>nx1002);
   ix4214 : mux21 port map ( Y=>nx4213, A0=>nx4215, A1=>nx4063, S0=>nx1012);
   ix1003 : xnor2 port map ( Y=>nx1002, A0=>nx4218, A1=>nx998);
   ix4219 : nand02 port map ( Y=>nx4218, A0=>nx5476, A1=>nx146);
   ix999 : xnor2 port map ( Y=>nx998, A0=>nx4221, A1=>nx770);
   ix4222 : mux21 port map ( Y=>nx4221, A0=>nx4223, A1=>nx4071, S0=>nx780);
   ix771 : xnor2 port map ( Y=>nx770, A0=>nx4227, A1=>nx766);
   ix4228 : nand02 port map ( Y=>nx4227, A0=>nx5472, A1=>nx122);
   ix767 : xnor2 port map ( Y=>nx766, A0=>nx4231, A1=>nx532);
   ix4232 : mux21 port map ( Y=>nx4231, A0=>nx4233, A1=>nx4077, S0=>nx548);
   ix533 : xnor2 port map ( Y=>nx532, A0=>nx4237, A1=>nx520);
   ix4240 : aoi22 port map ( Y=>nx4239, A0=>nx4022, A1=>mac_unit_tempP_16, 
      B0=>nx1911, B1=>nx4014);
   ix4443 : nor02ii port map ( Y=>mac_output(18), A0=>RST, A1=>nx4438);
   ix4439 : nor02 port map ( Y=>nx4438, A0=>RST, A1=>nx4251);
   ix4252 : xnor2 port map ( Y=>nx4251, A0=>nx4253, A1=>nx4257);
   ix4254 : xnor2 port map ( Y=>nx4253, A0=>mac_unit_tempP_18, A1=>nx4058);
   mac_unit_MR_reg_Q_18 : dffr port map ( Q=>mac_unit_tempP_18, QB=>OPEN, D
      =>nx4052, CLK=>CLK, R=>RST);
   ix4258 : mux21 port map ( Y=>nx4257, A0=>nx4105, A1=>nx4239, S0=>nx1909);
   ix4059 : xnor2 port map ( Y=>nx4058, A0=>nx4261, A1=>nx3544);
   ix4262 : mux21 port map ( Y=>nx4261, A0=>nx4107, A1=>nx4115, S0=>nx4111);
   ix3545 : xnor2 port map ( Y=>nx3544, A0=>nx4265, A1=>nx3540);
   ix4266 : nand02 port map ( Y=>nx4265, A0=>nx386, A1=>nx5520);
   ix3541 : xnor2 port map ( Y=>nx3540, A0=>nx3364, A1=>nx4271);
   ix3365 : mux21 port map ( Y=>nx3364, A0=>nx3318, A1=>nx3360, S0=>nx3322);
   ix4272 : xnor2 port map ( Y=>nx4271, A0=>nx4273, A1=>nx4275);
   ix4274 : nand02 port map ( Y=>nx4273, A0=>nx362, A1=>nx5516);
   ix4276 : xnor2 port map ( Y=>nx4275, A0=>nx4277, A1=>nx4281);
   ix4278 : mux21 port map ( Y=>nx4277, A0=>nx4279, A1=>nx4125, S0=>nx3090);
   ix4282 : xnor2 port map ( Y=>nx4281, A0=>nx4283, A1=>nx4285);
   ix4284 : nand02 port map ( Y=>nx4283, A0=>nx338, A1=>nx5512);
   ix4286 : xnor2 port map ( Y=>nx4285, A0=>nx4287, A1=>nx4291);
   ix4288 : mux21 port map ( Y=>nx4287, A0=>nx4289, A1=>nx4135, S0=>nx2858);
   ix4292 : xnor2 port map ( Y=>nx4291, A0=>nx4293, A1=>nx4295);
   ix4294 : nand02 port map ( Y=>nx4293, A0=>nx314, A1=>nx5508);
   ix4296 : xnor2 port map ( Y=>nx4295, A0=>nx4297, A1=>nx4301);
   ix4298 : mux21 port map ( Y=>nx4297, A0=>nx4299, A1=>nx4145, S0=>nx2626);
   ix4302 : xnor2 port map ( Y=>nx4301, A0=>nx4303, A1=>nx4305);
   ix4304 : nand02 port map ( Y=>nx4303, A0=>nx290, A1=>nx5504);
   ix4306 : xnor2 port map ( Y=>nx4305, A0=>nx4307, A1=>nx4311);
   ix4308 : mux21 port map ( Y=>nx4307, A0=>nx4309, A1=>nx4155, S0=>nx2394);
   ix4312 : xnor2 port map ( Y=>nx4311, A0=>nx4313, A1=>nx4315);
   ix4314 : nand02 port map ( Y=>nx4313, A0=>nx266, A1=>nx5500);
   ix4316 : xnor2 port map ( Y=>nx4315, A0=>nx4317, A1=>nx4321);
   ix4318 : mux21 port map ( Y=>nx4317, A0=>nx4319, A1=>nx4164, S0=>nx2162);
   ix4322 : xnor2 port map ( Y=>nx4321, A0=>nx4323, A1=>nx4325);
   ix4324 : nand02 port map ( Y=>nx4323, A0=>nx5496, A1=>nx242);
   ix4326 : xnor2 port map ( Y=>nx4325, A0=>nx4327, A1=>nx4331);
   ix4328 : mux21 port map ( Y=>nx4327, A0=>nx4329, A1=>nx4175, S0=>nx1930);
   ix4332 : xnor2 port map ( Y=>nx4331, A0=>nx4333, A1=>nx4335);
   ix4334 : nand02 port map ( Y=>nx4333, A0=>nx5492, A1=>nx218);
   ix4336 : xnor2 port map ( Y=>nx4335, A0=>nx4337, A1=>nx4341);
   ix4338 : mux21 port map ( Y=>nx4337, A0=>nx4339, A1=>nx4185, S0=>nx1698);
   ix4342 : xnor2 port map ( Y=>nx4341, A0=>nx4343, A1=>nx4345);
   ix4344 : nand02 port map ( Y=>nx4343, A0=>nx5488, A1=>nx194);
   ix4346 : xnor2 port map ( Y=>nx4345, A0=>nx4347, A1=>nx4351);
   ix4348 : mux21 port map ( Y=>nx4347, A0=>nx4349, A1=>nx4195, S0=>nx1466);
   ix4352 : xnor2 port map ( Y=>nx4351, A0=>nx4353, A1=>nx4355);
   ix4354 : nand02 port map ( Y=>nx4353, A0=>nx5484, A1=>nx170);
   ix4356 : xnor2 port map ( Y=>nx4355, A0=>nx4357, A1=>nx4361);
   ix4358 : mux21 port map ( Y=>nx4357, A0=>nx4359, A1=>nx4203, S0=>nx1234);
   ix4362 : xnor2 port map ( Y=>nx4361, A0=>nx4363, A1=>nx4365);
   ix4364 : nand02 port map ( Y=>nx4363, A0=>nx5480, A1=>nx146);
   ix4366 : xnor2 port map ( Y=>nx4365, A0=>nx4367, A1=>nx4371);
   ix4368 : mux21 port map ( Y=>nx4367, A0=>nx4369, A1=>nx4213, S0=>nx1002);
   ix4372 : xnor2 port map ( Y=>nx4371, A0=>nx4373, A1=>nx4375);
   ix4374 : nand02 port map ( Y=>nx4373, A0=>nx5476, A1=>nx122);
   ix4376 : xnor2 port map ( Y=>nx4375, A0=>nx4377, A1=>nx4381);
   ix4378 : mux21 port map ( Y=>nx4377, A0=>nx4379, A1=>nx4221, S0=>nx770);
   ix4382 : xnor2 port map ( Y=>nx4381, A0=>nx4383, A1=>nx4385);
   ix4386 : mux21 port map ( Y=>nx4385, A0=>nx4387, A1=>nx4231, S0=>nx532);
   ix4451 : nor02 port map ( Y=>mac_output(19), A0=>RST, A1=>nx4391);
   ix4392 : nand02 port map ( Y=>nx4391, A0=>nx2523, A1=>nx4070);
   ix4071 : xnor2 port map ( Y=>nx4070, A0=>nx1905, A1=>nx4501);
   ix4079 : xnor2 port map ( Y=>nx1905, A0=>mac_unit_tempP_19, A1=>nx4399);
   mac_unit_MR_reg_Q_19 : dffr port map ( Q=>mac_unit_tempP_19, QB=>OPEN, D
      =>nx4070, CLK=>CLK, R=>RST);
   ix4400 : xnor2 port map ( Y=>nx4399, A0=>nx4401, A1=>nx4405);
   ix4402 : mux21 port map ( Y=>nx4401, A0=>nx4403, A1=>nx4261, S0=>nx3544);
   ix4406 : xnor2 port map ( Y=>nx4405, A0=>nx4407, A1=>nx4409);
   ix4408 : nand02 port map ( Y=>nx4407, A0=>nx362, A1=>nx5520);
   ix4410 : xnor2 port map ( Y=>nx4409, A0=>nx4411, A1=>nx4415);
   ix4412 : mux21 port map ( Y=>nx4411, A0=>nx4413, A1=>nx4275, S0=>nx4271);
   ix4416 : xnor2 port map ( Y=>nx4415, A0=>nx4417, A1=>nx4419);
   ix4418 : nand02 port map ( Y=>nx4417, A0=>nx338, A1=>nx5516);
   ix4420 : xnor2 port map ( Y=>nx4419, A0=>nx4421, A1=>nx4423);
   ix4422 : mux21 port map ( Y=>nx4421, A0=>nx4277, A1=>nx4285, S0=>nx4281);
   ix4424 : xnor2 port map ( Y=>nx4423, A0=>nx4425, A1=>nx4427);
   ix4426 : nand02 port map ( Y=>nx4425, A0=>nx314, A1=>nx5512);
   ix4428 : xnor2 port map ( Y=>nx4427, A0=>nx4429, A1=>nx4431);
   ix4430 : mux21 port map ( Y=>nx4429, A0=>nx4287, A1=>nx4295, S0=>nx4291);
   ix4432 : xnor2 port map ( Y=>nx4431, A0=>nx4433, A1=>nx4435);
   ix4434 : nand02 port map ( Y=>nx4433, A0=>nx290, A1=>nx5508);
   ix4436 : xnor2 port map ( Y=>nx4435, A0=>nx4437, A1=>nx4439);
   ix4438 : mux21 port map ( Y=>nx4437, A0=>nx4297, A1=>nx4305, S0=>nx4301);
   ix4440 : xnor2 port map ( Y=>nx4439, A0=>nx4441, A1=>nx4443);
   ix4442 : nand02 port map ( Y=>nx4441, A0=>nx266, A1=>nx5504);
   ix4444 : xnor2 port map ( Y=>nx4443, A0=>nx4445, A1=>nx4447);
   ix4446 : mux21 port map ( Y=>nx4445, A0=>nx4307, A1=>nx4315, S0=>nx4311);
   ix4448 : xnor2 port map ( Y=>nx4447, A0=>nx4449, A1=>nx4451);
   ix4450 : nand02 port map ( Y=>nx4449, A0=>nx242, A1=>nx5500);
   ix4452 : xnor2 port map ( Y=>nx4451, A0=>nx4453, A1=>nx4455);
   ix4454 : mux21 port map ( Y=>nx4453, A0=>nx4317, A1=>nx4325, S0=>nx4321);
   ix4456 : xnor2 port map ( Y=>nx4455, A0=>nx4457, A1=>nx4459);
   ix4458 : nand02 port map ( Y=>nx4457, A0=>nx5496, A1=>nx218);
   ix4460 : xnor2 port map ( Y=>nx4459, A0=>nx4461, A1=>nx4463);
   ix4462 : mux21 port map ( Y=>nx4461, A0=>nx4327, A1=>nx4335, S0=>nx4331);
   ix4464 : xnor2 port map ( Y=>nx4463, A0=>nx4465, A1=>nx4467);
   ix4466 : nand02 port map ( Y=>nx4465, A0=>nx5492, A1=>nx194);
   ix4468 : xnor2 port map ( Y=>nx4467, A0=>nx4469, A1=>nx4471);
   ix4470 : mux21 port map ( Y=>nx4469, A0=>nx4337, A1=>nx4345, S0=>nx4341);
   ix4472 : xnor2 port map ( Y=>nx4471, A0=>nx4473, A1=>nx4475);
   ix4474 : nand02 port map ( Y=>nx4473, A0=>nx5488, A1=>nx170);
   ix4476 : xnor2 port map ( Y=>nx4475, A0=>nx4477, A1=>nx4479);
   ix4478 : mux21 port map ( Y=>nx4477, A0=>nx4347, A1=>nx4355, S0=>nx4351);
   ix4480 : xnor2 port map ( Y=>nx4479, A0=>nx4481, A1=>nx4483);
   ix4482 : nand02 port map ( Y=>nx4481, A0=>nx5484, A1=>nx146);
   ix4484 : xnor2 port map ( Y=>nx4483, A0=>nx4485, A1=>nx4487);
   ix4486 : mux21 port map ( Y=>nx4485, A0=>nx4357, A1=>nx4365, S0=>nx4361);
   ix4488 : xnor2 port map ( Y=>nx4487, A0=>nx4489, A1=>nx4491);
   ix4490 : nand02 port map ( Y=>nx4489, A0=>nx5480, A1=>nx122);
   ix4492 : xnor2 port map ( Y=>nx4491, A0=>nx4493, A1=>nx4495);
   ix4494 : mux21 port map ( Y=>nx4493, A0=>nx4367, A1=>nx4375, S0=>nx4371);
   ix4496 : xnor2 port map ( Y=>nx4495, A0=>nx4497, A1=>nx4499);
   ix4500 : mux21 port map ( Y=>nx4499, A0=>nx4377, A1=>nx4385, S0=>nx4381);
   ix4502 : aoi22 port map ( Y=>nx4501, A0=>nx4058, A1=>mac_unit_tempP_18, 
      B0=>nx1907, B1=>nx4050);
   ix4459 : nor02 port map ( Y=>mac_output(20), A0=>RST, A1=>nx4511);
   ix4512 : nand02 port map ( Y=>nx4511, A0=>nx2523, A1=>nx4088);
   ix4089 : xnor2 port map ( Y=>nx4088, A0=>nx1903, A1=>nx4609);
   ix4097 : xnor2 port map ( Y=>nx1903, A0=>mac_unit_tempP_20, A1=>nx4519);
   mac_unit_MR_reg_Q_20 : dffr port map ( Q=>mac_unit_tempP_20, QB=>OPEN, D
      =>nx4088, CLK=>CLK, R=>RST);
   ix4520 : xnor2 port map ( Y=>nx4519, A0=>nx4521, A1=>nx4523);
   ix4522 : mux21 port map ( Y=>nx4521, A0=>nx4401, A1=>nx4409, S0=>nx4405);
   ix4524 : xnor2 port map ( Y=>nx4523, A0=>nx4525, A1=>nx4527);
   ix4526 : nand02 port map ( Y=>nx4525, A0=>nx338, A1=>nx5520);
   ix4528 : xnor2 port map ( Y=>nx4527, A0=>nx4529, A1=>nx4531);
   ix4530 : mux21 port map ( Y=>nx4529, A0=>nx4411, A1=>nx4419, S0=>nx4415);
   ix4532 : xnor2 port map ( Y=>nx4531, A0=>nx4533, A1=>nx4535);
   ix4534 : nand02 port map ( Y=>nx4533, A0=>nx314, A1=>nx5516);
   ix4536 : xnor2 port map ( Y=>nx4535, A0=>nx4537, A1=>nx4539);
   ix4538 : mux21 port map ( Y=>nx4537, A0=>nx4421, A1=>nx4427, S0=>nx4423);
   ix4540 : xnor2 port map ( Y=>nx4539, A0=>nx4541, A1=>nx4543);
   ix4542 : nand02 port map ( Y=>nx4541, A0=>nx290, A1=>nx5512);
   ix4544 : xnor2 port map ( Y=>nx4543, A0=>nx4545, A1=>nx4547);
   ix4546 : mux21 port map ( Y=>nx4545, A0=>nx4429, A1=>nx4435, S0=>nx4431);
   ix4548 : xnor2 port map ( Y=>nx4547, A0=>nx4549, A1=>nx4551);
   ix4550 : nand02 port map ( Y=>nx4549, A0=>nx266, A1=>nx5508);
   ix4552 : xnor2 port map ( Y=>nx4551, A0=>nx4553, A1=>nx4555);
   ix4554 : mux21 port map ( Y=>nx4553, A0=>nx4437, A1=>nx4443, S0=>nx4439);
   ix4556 : xnor2 port map ( Y=>nx4555, A0=>nx4557, A1=>nx4559);
   ix4558 : nand02 port map ( Y=>nx4557, A0=>nx242, A1=>nx5504);
   ix4560 : xnor2 port map ( Y=>nx4559, A0=>nx4561, A1=>nx4563);
   ix4562 : mux21 port map ( Y=>nx4561, A0=>nx4445, A1=>nx4451, S0=>nx4447);
   ix4564 : xnor2 port map ( Y=>nx4563, A0=>nx4565, A1=>nx4567);
   ix4566 : nand02 port map ( Y=>nx4565, A0=>nx5500, A1=>nx218);
   ix4568 : xnor2 port map ( Y=>nx4567, A0=>nx4569, A1=>nx4571);
   ix4570 : mux21 port map ( Y=>nx4569, A0=>nx4453, A1=>nx4459, S0=>nx4455);
   ix4572 : xnor2 port map ( Y=>nx4571, A0=>nx4573, A1=>nx4575);
   ix4574 : nand02 port map ( Y=>nx4573, A0=>nx5496, A1=>nx194);
   ix4576 : xnor2 port map ( Y=>nx4575, A0=>nx4577, A1=>nx4579);
   ix4578 : mux21 port map ( Y=>nx4577, A0=>nx4461, A1=>nx4467, S0=>nx4463);
   ix4580 : xnor2 port map ( Y=>nx4579, A0=>nx4581, A1=>nx4583);
   ix4582 : nand02 port map ( Y=>nx4581, A0=>nx5492, A1=>nx170);
   ix4584 : xnor2 port map ( Y=>nx4583, A0=>nx4585, A1=>nx4587);
   ix4586 : mux21 port map ( Y=>nx4585, A0=>nx4469, A1=>nx4475, S0=>nx4471);
   ix4588 : xnor2 port map ( Y=>nx4587, A0=>nx4589, A1=>nx4591);
   ix4590 : nand02 port map ( Y=>nx4589, A0=>nx5488, A1=>nx146);
   ix4592 : xnor2 port map ( Y=>nx4591, A0=>nx4593, A1=>nx4595);
   ix4594 : mux21 port map ( Y=>nx4593, A0=>nx4477, A1=>nx4483, S0=>nx4479);
   ix4596 : xnor2 port map ( Y=>nx4595, A0=>nx4597, A1=>nx4599);
   ix4598 : nand02 port map ( Y=>nx4597, A0=>nx5484, A1=>nx122);
   ix4600 : xnor2 port map ( Y=>nx4599, A0=>nx4601, A1=>nx4603);
   ix4602 : mux21 port map ( Y=>nx4601, A0=>nx4485, A1=>nx4491, S0=>nx4487);
   ix4604 : xnor2 port map ( Y=>nx4603, A0=>nx4605, A1=>nx4607);
   ix4608 : mux21 port map ( Y=>nx4607, A0=>nx4493, A1=>nx4499, S0=>nx4495);
   ix4610 : mux21 port map ( Y=>nx4609, A0=>nx4399, A1=>nx4501, S0=>nx1905);
   ix4467 : nor02 port map ( Y=>mac_output(21), A0=>RST, A1=>nx4613);
   ix4614 : nand02 port map ( Y=>nx4613, A0=>nx2523, A1=>nx4106);
   ix4107 : xnor2 port map ( Y=>nx4106, A0=>nx1902, A1=>nx4703);
   ix4115 : xnor2 port map ( Y=>nx1902, A0=>mac_unit_tempP_21, A1=>nx4620);
   mac_unit_MR_reg_Q_21 : dffr port map ( Q=>mac_unit_tempP_21, QB=>OPEN, D
      =>nx4106, CLK=>CLK, R=>RST);
   ix4621 : xnor2 port map ( Y=>nx4620, A0=>nx4623, A1=>nx4625);
   ix4624 : mux21 port map ( Y=>nx4623, A0=>nx4521, A1=>nx4527, S0=>nx4523);
   ix4626 : xnor2 port map ( Y=>nx4625, A0=>nx4627, A1=>nx4629);
   ix4628 : nand02 port map ( Y=>nx4627, A0=>nx314, A1=>nx5520);
   ix4630 : xnor2 port map ( Y=>nx4629, A0=>nx4631, A1=>nx4633);
   ix4632 : mux21 port map ( Y=>nx4631, A0=>nx4529, A1=>nx4535, S0=>nx4531);
   ix4634 : xnor2 port map ( Y=>nx4633, A0=>nx4635, A1=>nx4637);
   ix4636 : nand02 port map ( Y=>nx4635, A0=>nx290, A1=>nx5516);
   ix4638 : xnor2 port map ( Y=>nx4637, A0=>nx4639, A1=>nx4641);
   ix4640 : mux21 port map ( Y=>nx4639, A0=>nx4537, A1=>nx4543, S0=>nx4539);
   ix4642 : xnor2 port map ( Y=>nx4641, A0=>nx4643, A1=>nx4645);
   ix4644 : nand02 port map ( Y=>nx4643, A0=>nx266, A1=>nx5512);
   ix4646 : xnor2 port map ( Y=>nx4645, A0=>nx4647, A1=>nx4649);
   ix4648 : mux21 port map ( Y=>nx4647, A0=>nx4545, A1=>nx4551, S0=>nx4547);
   ix4650 : xnor2 port map ( Y=>nx4649, A0=>nx4651, A1=>nx4653);
   ix4652 : nand02 port map ( Y=>nx4651, A0=>nx242, A1=>nx5508);
   ix4654 : xnor2 port map ( Y=>nx4653, A0=>nx4655, A1=>nx4657);
   ix4656 : mux21 port map ( Y=>nx4655, A0=>nx4553, A1=>nx4559, S0=>nx4555);
   ix4658 : xnor2 port map ( Y=>nx4657, A0=>nx4659, A1=>nx4661);
   ix4660 : nand02 port map ( Y=>nx4659, A0=>nx218, A1=>nx5504);
   ix4662 : xnor2 port map ( Y=>nx4661, A0=>nx4663, A1=>nx4665);
   ix4664 : mux21 port map ( Y=>nx4663, A0=>nx4561, A1=>nx4567, S0=>nx4563);
   ix4666 : xnor2 port map ( Y=>nx4665, A0=>nx4667, A1=>nx4669);
   ix4668 : nand02 port map ( Y=>nx4667, A0=>nx5500, A1=>nx194);
   ix4670 : xnor2 port map ( Y=>nx4669, A0=>nx4671, A1=>nx4673);
   ix4672 : mux21 port map ( Y=>nx4671, A0=>nx4569, A1=>nx4575, S0=>nx4571);
   ix4674 : xnor2 port map ( Y=>nx4673, A0=>nx4675, A1=>nx4677);
   ix4676 : nand02 port map ( Y=>nx4675, A0=>nx5496, A1=>nx170);
   ix4678 : xnor2 port map ( Y=>nx4677, A0=>nx4679, A1=>nx4681);
   ix4680 : mux21 port map ( Y=>nx4679, A0=>nx4577, A1=>nx4583, S0=>nx4579);
   ix4682 : xnor2 port map ( Y=>nx4681, A0=>nx4683, A1=>nx4685);
   ix4684 : nand02 port map ( Y=>nx4683, A0=>nx5492, A1=>nx146);
   ix4686 : xnor2 port map ( Y=>nx4685, A0=>nx4687, A1=>nx4689);
   ix4688 : mux21 port map ( Y=>nx4687, A0=>nx4585, A1=>nx4591, S0=>nx4587);
   ix4690 : xnor2 port map ( Y=>nx4689, A0=>nx4691, A1=>nx4693);
   ix4692 : nand02 port map ( Y=>nx4691, A0=>nx5488, A1=>nx122);
   ix4694 : xnor2 port map ( Y=>nx4693, A0=>nx4695, A1=>nx4697);
   ix4696 : mux21 port map ( Y=>nx4695, A0=>nx4593, A1=>nx4599, S0=>nx4595);
   ix4698 : xnor2 port map ( Y=>nx4697, A0=>nx4699, A1=>nx4701);
   ix4702 : mux21 port map ( Y=>nx4701, A0=>nx4601, A1=>nx4607, S0=>nx4603);
   ix4704 : mux21 port map ( Y=>nx4703, A0=>nx4519, A1=>nx4609, S0=>nx1903);
   ix4475 : nor02 port map ( Y=>mac_output(22), A0=>RST, A1=>nx4707);
   ix4708 : nand02 port map ( Y=>nx4707, A0=>nx2523, A1=>nx4124);
   ix4125 : xnor2 port map ( Y=>nx4124, A0=>nx1901, A1=>nx4789);
   ix4133 : xnor2 port map ( Y=>nx1901, A0=>mac_unit_tempP_22, A1=>nx4714);
   mac_unit_MR_reg_Q_22 : dffr port map ( Q=>mac_unit_tempP_22, QB=>OPEN, D
      =>nx4124, CLK=>CLK, R=>RST);
   ix4715 : xnor2 port map ( Y=>nx4714, A0=>nx4716, A1=>nx4719);
   ix4717 : mux21 port map ( Y=>nx4716, A0=>nx4623, A1=>nx4629, S0=>nx4625);
   ix4720 : xnor2 port map ( Y=>nx4719, A0=>nx4721, A1=>nx4723);
   ix4722 : nand02 port map ( Y=>nx4721, A0=>nx290, A1=>nx5520);
   ix4724 : xnor2 port map ( Y=>nx4723, A0=>nx4725, A1=>nx4727);
   ix4726 : mux21 port map ( Y=>nx4725, A0=>nx4631, A1=>nx4637, S0=>nx4633);
   ix4728 : xnor2 port map ( Y=>nx4727, A0=>nx4729, A1=>nx4731);
   ix4730 : nand02 port map ( Y=>nx4729, A0=>nx266, A1=>nx5516);
   ix4732 : xnor2 port map ( Y=>nx4731, A0=>nx4733, A1=>nx4735);
   ix4734 : mux21 port map ( Y=>nx4733, A0=>nx4639, A1=>nx4645, S0=>nx4641);
   ix4736 : xnor2 port map ( Y=>nx4735, A0=>nx4737, A1=>nx4739);
   ix4738 : nand02 port map ( Y=>nx4737, A0=>nx242, A1=>nx5512);
   ix4740 : xnor2 port map ( Y=>nx4739, A0=>nx4741, A1=>nx4743);
   ix4742 : mux21 port map ( Y=>nx4741, A0=>nx4647, A1=>nx4653, S0=>nx4649);
   ix4744 : xnor2 port map ( Y=>nx4743, A0=>nx4745, A1=>nx4747);
   ix4746 : nand02 port map ( Y=>nx4745, A0=>nx218, A1=>nx5508);
   ix4748 : xnor2 port map ( Y=>nx4747, A0=>nx4749, A1=>nx4751);
   ix4750 : mux21 port map ( Y=>nx4749, A0=>nx4655, A1=>nx4661, S0=>nx4657);
   ix4752 : xnor2 port map ( Y=>nx4751, A0=>nx4753, A1=>nx4755);
   ix4754 : nand02 port map ( Y=>nx4753, A0=>nx5504, A1=>nx194);
   ix4756 : xnor2 port map ( Y=>nx4755, A0=>nx4757, A1=>nx4759);
   ix4758 : mux21 port map ( Y=>nx4757, A0=>nx4663, A1=>nx4669, S0=>nx4665);
   ix4760 : xnor2 port map ( Y=>nx4759, A0=>nx4761, A1=>nx4763);
   ix4762 : nand02 port map ( Y=>nx4761, A0=>nx5500, A1=>nx170);
   ix4764 : xnor2 port map ( Y=>nx4763, A0=>nx4765, A1=>nx4767);
   ix4766 : mux21 port map ( Y=>nx4765, A0=>nx4671, A1=>nx4677, S0=>nx4673);
   ix4768 : xnor2 port map ( Y=>nx4767, A0=>nx4769, A1=>nx4771);
   ix4770 : nand02 port map ( Y=>nx4769, A0=>nx5496, A1=>nx146);
   ix4772 : xnor2 port map ( Y=>nx4771, A0=>nx4773, A1=>nx4775);
   ix4774 : mux21 port map ( Y=>nx4773, A0=>nx4679, A1=>nx4685, S0=>nx4681);
   ix4776 : xnor2 port map ( Y=>nx4775, A0=>nx4777, A1=>nx4779);
   ix4778 : nand02 port map ( Y=>nx4777, A0=>nx5492, A1=>nx122);
   ix4780 : xnor2 port map ( Y=>nx4779, A0=>nx4781, A1=>nx4783);
   ix4782 : mux21 port map ( Y=>nx4781, A0=>nx4687, A1=>nx4693, S0=>nx4689);
   ix4784 : xnor2 port map ( Y=>nx4783, A0=>nx4785, A1=>nx4787);
   ix4788 : mux21 port map ( Y=>nx4787, A0=>nx4695, A1=>nx4701, S0=>nx4697);
   ix4790 : mux21 port map ( Y=>nx4789, A0=>nx4620, A1=>nx4703, S0=>nx1902);
   ix4483 : nor02 port map ( Y=>mac_output(23), A0=>RST, A1=>nx4793);
   ix4794 : nand02 port map ( Y=>nx4793, A0=>nx2523, A1=>nx4142);
   ix4143 : xnor2 port map ( Y=>nx4142, A0=>nx1899, A1=>nx4865);
   ix4151 : xnor2 port map ( Y=>nx1899, A0=>mac_unit_tempP_23, A1=>nx4799);
   mac_unit_MR_reg_Q_23 : dffr port map ( Q=>mac_unit_tempP_23, QB=>OPEN, D
      =>nx4142, CLK=>CLK, R=>RST);
   ix4800 : xnor2 port map ( Y=>nx4799, A0=>nx4801, A1=>nx4803);
   ix4802 : mux21 port map ( Y=>nx4801, A0=>nx4716, A1=>nx4723, S0=>nx4719);
   ix4804 : xnor2 port map ( Y=>nx4803, A0=>nx4805, A1=>nx4807);
   ix4806 : nand02 port map ( Y=>nx4805, A0=>nx266, A1=>nx5520);
   ix4808 : xnor2 port map ( Y=>nx4807, A0=>nx4809, A1=>nx4811);
   ix4810 : mux21 port map ( Y=>nx4809, A0=>nx4725, A1=>nx4731, S0=>nx4727);
   ix4812 : xnor2 port map ( Y=>nx4811, A0=>nx4813, A1=>nx4815);
   ix4814 : nand02 port map ( Y=>nx4813, A0=>nx242, A1=>nx5516);
   ix4816 : xnor2 port map ( Y=>nx4815, A0=>nx4817, A1=>nx4819);
   ix4818 : mux21 port map ( Y=>nx4817, A0=>nx4733, A1=>nx4739, S0=>nx4735);
   ix4820 : xnor2 port map ( Y=>nx4819, A0=>nx4821, A1=>nx4823);
   ix4822 : nand02 port map ( Y=>nx4821, A0=>nx218, A1=>nx5512);
   ix4824 : xnor2 port map ( Y=>nx4823, A0=>nx4825, A1=>nx4827);
   ix4826 : mux21 port map ( Y=>nx4825, A0=>nx4741, A1=>nx4747, S0=>nx4743);
   ix4828 : xnor2 port map ( Y=>nx4827, A0=>nx4829, A1=>nx4831);
   ix4830 : nand02 port map ( Y=>nx4829, A0=>nx194, A1=>nx5508);
   ix4832 : xnor2 port map ( Y=>nx4831, A0=>nx4833, A1=>nx4835);
   ix4834 : mux21 port map ( Y=>nx4833, A0=>nx4749, A1=>nx4755, S0=>nx4751);
   ix4836 : xnor2 port map ( Y=>nx4835, A0=>nx4837, A1=>nx4839);
   ix4838 : nand02 port map ( Y=>nx4837, A0=>nx5504, A1=>nx170);
   ix4840 : xnor2 port map ( Y=>nx4839, A0=>nx4841, A1=>nx4843);
   ix4842 : mux21 port map ( Y=>nx4841, A0=>nx4757, A1=>nx4763, S0=>nx4759);
   ix4844 : xnor2 port map ( Y=>nx4843, A0=>nx4845, A1=>nx4847);
   ix4846 : nand02 port map ( Y=>nx4845, A0=>nx5500, A1=>nx146);
   ix4848 : xnor2 port map ( Y=>nx4847, A0=>nx4849, A1=>nx4851);
   ix4850 : mux21 port map ( Y=>nx4849, A0=>nx4765, A1=>nx4771, S0=>nx4767);
   ix4852 : xnor2 port map ( Y=>nx4851, A0=>nx4853, A1=>nx4855);
   ix4854 : nand02 port map ( Y=>nx4853, A0=>nx5496, A1=>nx122);
   ix4856 : xnor2 port map ( Y=>nx4855, A0=>nx4857, A1=>nx4859);
   ix4858 : mux21 port map ( Y=>nx4857, A0=>nx4773, A1=>nx4779, S0=>nx4775);
   ix4860 : xnor2 port map ( Y=>nx4859, A0=>nx4861, A1=>nx4863);
   ix4864 : mux21 port map ( Y=>nx4863, A0=>nx4781, A1=>nx4787, S0=>nx4783);
   ix4866 : mux21 port map ( Y=>nx4865, A0=>nx4714, A1=>nx4789, S0=>nx1901);
   ix4491 : nor02 port map ( Y=>mac_output(24), A0=>RST, A1=>nx4868);
   ix4869 : nand02 port map ( Y=>nx4868, A0=>nx2523, A1=>nx4160);
   ix4161 : xnor2 port map ( Y=>nx4160, A0=>nx1897, A1=>nx4933);
   ix4169 : xnor2 port map ( Y=>nx1897, A0=>mac_unit_tempP_24, A1=>nx4875);
   mac_unit_MR_reg_Q_24 : dffr port map ( Q=>mac_unit_tempP_24, QB=>OPEN, D
      =>nx4160, CLK=>CLK, R=>RST);
   ix4876 : xnor2 port map ( Y=>nx4875, A0=>nx4877, A1=>nx4879);
   ix4878 : mux21 port map ( Y=>nx4877, A0=>nx4801, A1=>nx4807, S0=>nx4803);
   ix4880 : xnor2 port map ( Y=>nx4879, A0=>nx4881, A1=>nx4883);
   ix4882 : nand02 port map ( Y=>nx4881, A0=>nx242, A1=>nx5520);
   ix4884 : xnor2 port map ( Y=>nx4883, A0=>nx4885, A1=>nx4887);
   ix4886 : mux21 port map ( Y=>nx4885, A0=>nx4809, A1=>nx4815, S0=>nx4811);
   ix4888 : xnor2 port map ( Y=>nx4887, A0=>nx4889, A1=>nx4891);
   ix4890 : nand02 port map ( Y=>nx4889, A0=>nx218, A1=>nx5516);
   ix4892 : xnor2 port map ( Y=>nx4891, A0=>nx4893, A1=>nx4895);
   ix4894 : mux21 port map ( Y=>nx4893, A0=>nx4817, A1=>nx4823, S0=>nx4819);
   ix4896 : xnor2 port map ( Y=>nx4895, A0=>nx4897, A1=>nx4899);
   ix4898 : nand02 port map ( Y=>nx4897, A0=>nx194, A1=>nx5512);
   ix4900 : xnor2 port map ( Y=>nx4899, A0=>nx4901, A1=>nx4903);
   ix4902 : mux21 port map ( Y=>nx4901, A0=>nx4825, A1=>nx4831, S0=>nx4827);
   ix4904 : xnor2 port map ( Y=>nx4903, A0=>nx4905, A1=>nx4907);
   ix4906 : nand02 port map ( Y=>nx4905, A0=>nx5508, A1=>nx170);
   ix4908 : xnor2 port map ( Y=>nx4907, A0=>nx4909, A1=>nx4911);
   ix4910 : mux21 port map ( Y=>nx4909, A0=>nx4833, A1=>nx4839, S0=>nx4835);
   ix4912 : xnor2 port map ( Y=>nx4911, A0=>nx4913, A1=>nx4915);
   ix4914 : nand02 port map ( Y=>nx4913, A0=>nx5504, A1=>nx146);
   ix4916 : xnor2 port map ( Y=>nx4915, A0=>nx4917, A1=>nx4919);
   ix4918 : mux21 port map ( Y=>nx4917, A0=>nx4841, A1=>nx4847, S0=>nx4843);
   ix4920 : xnor2 port map ( Y=>nx4919, A0=>nx4921, A1=>nx4923);
   ix4922 : nand02 port map ( Y=>nx4921, A0=>nx5500, A1=>nx122);
   ix4924 : xnor2 port map ( Y=>nx4923, A0=>nx4925, A1=>nx4927);
   ix4926 : mux21 port map ( Y=>nx4925, A0=>nx4849, A1=>nx4855, S0=>nx4851);
   ix4928 : xnor2 port map ( Y=>nx4927, A0=>nx4929, A1=>nx4931);
   ix4932 : mux21 port map ( Y=>nx4931, A0=>nx4857, A1=>nx4863, S0=>nx4859);
   ix4934 : mux21 port map ( Y=>nx4933, A0=>nx4799, A1=>nx4865, S0=>nx1899);
   ix4499 : nor02 port map ( Y=>mac_output(25), A0=>RST, A1=>nx4937);
   ix4938 : nand02 port map ( Y=>nx4937, A0=>nx2523, A1=>nx4178);
   ix4179 : xnor2 port map ( Y=>nx4178, A0=>nx1895, A1=>nx4993);
   ix4187 : xnor2 port map ( Y=>nx1895, A0=>mac_unit_tempP_25, A1=>nx4943);
   mac_unit_MR_reg_Q_25 : dffr port map ( Q=>mac_unit_tempP_25, QB=>OPEN, D
      =>nx4178, CLK=>CLK, R=>RST);
   ix4944 : xnor2 port map ( Y=>nx4943, A0=>nx4945, A1=>nx4947);
   ix4946 : mux21 port map ( Y=>nx4945, A0=>nx4877, A1=>nx4883, S0=>nx4879);
   ix4948 : xnor2 port map ( Y=>nx4947, A0=>nx4949, A1=>nx4951);
   ix4950 : nand02 port map ( Y=>nx4949, A0=>nx218, A1=>nx5520);
   ix4952 : xnor2 port map ( Y=>nx4951, A0=>nx4953, A1=>nx4955);
   ix4954 : mux21 port map ( Y=>nx4953, A0=>nx4885, A1=>nx4891, S0=>nx4887);
   ix4956 : xnor2 port map ( Y=>nx4955, A0=>nx4957, A1=>nx4959);
   ix4958 : nand02 port map ( Y=>nx4957, A0=>nx194, A1=>nx5516);
   ix4960 : xnor2 port map ( Y=>nx4959, A0=>nx4961, A1=>nx4963);
   ix4962 : mux21 port map ( Y=>nx4961, A0=>nx4893, A1=>nx4899, S0=>nx4895);
   ix4964 : xnor2 port map ( Y=>nx4963, A0=>nx4965, A1=>nx4967);
   ix4966 : nand02 port map ( Y=>nx4965, A0=>nx170, A1=>nx5512);
   ix4968 : xnor2 port map ( Y=>nx4967, A0=>nx4969, A1=>nx4971);
   ix4970 : mux21 port map ( Y=>nx4969, A0=>nx4901, A1=>nx4907, S0=>nx4903);
   ix4972 : xnor2 port map ( Y=>nx4971, A0=>nx4973, A1=>nx4975);
   ix4974 : nand02 port map ( Y=>nx4973, A0=>nx5508, A1=>nx146);
   ix4976 : xnor2 port map ( Y=>nx4975, A0=>nx4977, A1=>nx4979);
   ix4978 : mux21 port map ( Y=>nx4977, A0=>nx4909, A1=>nx4915, S0=>nx4911);
   ix4980 : xnor2 port map ( Y=>nx4979, A0=>nx4981, A1=>nx4983);
   ix4982 : nand02 port map ( Y=>nx4981, A0=>nx5504, A1=>nx122);
   ix4984 : xnor2 port map ( Y=>nx4983, A0=>nx4985, A1=>nx4987);
   ix4986 : mux21 port map ( Y=>nx4985, A0=>nx4917, A1=>nx4923, S0=>nx4919);
   ix4988 : xnor2 port map ( Y=>nx4987, A0=>nx4989, A1=>nx4991);
   ix4992 : mux21 port map ( Y=>nx4991, A0=>nx4925, A1=>nx4931, S0=>nx4927);
   ix4994 : mux21 port map ( Y=>nx4993, A0=>nx4875, A1=>nx4933, S0=>nx1897);
   ix4507 : nor02 port map ( Y=>mac_output(26), A0=>RST, A1=>nx4996);
   ix4997 : nand02 port map ( Y=>nx4996, A0=>nx2523, A1=>nx4196);
   ix4197 : xnor2 port map ( Y=>nx4196, A0=>nx1893, A1=>nx5044);
   ix4205 : xnor2 port map ( Y=>nx1893, A0=>mac_unit_tempP_26, A1=>nx5002);
   mac_unit_MR_reg_Q_26 : dffr port map ( Q=>mac_unit_tempP_26, QB=>OPEN, D
      =>nx4196, CLK=>CLK, R=>RST);
   ix5003 : xnor2 port map ( Y=>nx5002, A0=>nx5004, A1=>nx5006);
   ix5005 : mux21 port map ( Y=>nx5004, A0=>nx4945, A1=>nx4951, S0=>nx4947);
   ix5007 : xnor2 port map ( Y=>nx5006, A0=>nx5008, A1=>nx5010);
   ix5009 : nand02 port map ( Y=>nx5008, A0=>nx194, A1=>nx5520);
   ix5011 : xnor2 port map ( Y=>nx5010, A0=>nx5012, A1=>nx5014);
   ix5013 : mux21 port map ( Y=>nx5012, A0=>nx4953, A1=>nx4959, S0=>nx4955);
   ix5015 : xnor2 port map ( Y=>nx5014, A0=>nx5016, A1=>nx5018);
   ix5017 : nand02 port map ( Y=>nx5016, A0=>nx170, A1=>nx5516);
   ix5019 : xnor2 port map ( Y=>nx5018, A0=>nx5020, A1=>nx5022);
   ix5021 : mux21 port map ( Y=>nx5020, A0=>nx4961, A1=>nx4967, S0=>nx4963);
   ix5023 : xnor2 port map ( Y=>nx5022, A0=>nx5024, A1=>nx5026);
   ix5025 : nand02 port map ( Y=>nx5024, A0=>nx5512, A1=>nx146);
   ix5027 : xnor2 port map ( Y=>nx5026, A0=>nx5028, A1=>nx5030);
   ix5029 : mux21 port map ( Y=>nx5028, A0=>nx4969, A1=>nx4975, S0=>nx4971);
   ix5031 : xnor2 port map ( Y=>nx5030, A0=>nx5032, A1=>nx5034);
   ix5033 : nand02 port map ( Y=>nx5032, A0=>nx5508, A1=>nx122);
   ix5035 : xnor2 port map ( Y=>nx5034, A0=>nx5036, A1=>nx5038);
   ix5037 : mux21 port map ( Y=>nx5036, A0=>nx4977, A1=>nx4983, S0=>nx4979);
   ix5039 : xnor2 port map ( Y=>nx5038, A0=>nx5040, A1=>nx5042);
   ix5043 : mux21 port map ( Y=>nx5042, A0=>nx4985, A1=>nx4991, S0=>nx4987);
   ix5045 : mux21 port map ( Y=>nx5044, A0=>nx4943, A1=>nx4993, S0=>nx1895);
   ix4515 : nor02 port map ( Y=>mac_output(27), A0=>RST, A1=>nx5047);
   ix5048 : nand02 port map ( Y=>nx5047, A0=>nx2523, A1=>nx4214);
   ix4215 : xnor2 port map ( Y=>nx4214, A0=>nx1892, A1=>nx5087);
   ix4223 : xnor2 port map ( Y=>nx1892, A0=>mac_unit_tempP_27, A1=>nx5053);
   mac_unit_MR_reg_Q_27 : dffr port map ( Q=>mac_unit_tempP_27, QB=>OPEN, D
      =>nx4214, CLK=>CLK, R=>RST);
   ix5054 : xnor2 port map ( Y=>nx5053, A0=>nx5055, A1=>nx5057);
   ix5056 : mux21 port map ( Y=>nx5055, A0=>nx5004, A1=>nx5010, S0=>nx5006);
   ix5058 : xnor2 port map ( Y=>nx5057, A0=>nx5059, A1=>nx5061);
   ix5060 : nand02 port map ( Y=>nx5059, A0=>nx170, A1=>nx5520);
   ix5062 : xnor2 port map ( Y=>nx5061, A0=>nx5063, A1=>nx5065);
   ix5064 : mux21 port map ( Y=>nx5063, A0=>nx5012, A1=>nx5018, S0=>nx5014);
   ix5066 : xnor2 port map ( Y=>nx5065, A0=>nx5067, A1=>nx5069);
   ix5068 : nand02 port map ( Y=>nx5067, A0=>nx146, A1=>nx5516);
   ix5070 : xnor2 port map ( Y=>nx5069, A0=>nx5071, A1=>nx5073);
   ix5072 : mux21 port map ( Y=>nx5071, A0=>nx5020, A1=>nx5026, S0=>nx5022);
   ix5074 : xnor2 port map ( Y=>nx5073, A0=>nx5075, A1=>nx5077);
   ix5076 : nand02 port map ( Y=>nx5075, A0=>nx5512, A1=>nx122);
   ix5078 : xnor2 port map ( Y=>nx5077, A0=>nx5079, A1=>nx5081);
   ix5080 : mux21 port map ( Y=>nx5079, A0=>nx5028, A1=>nx5034, S0=>nx5030);
   ix5082 : xnor2 port map ( Y=>nx5081, A0=>nx5083, A1=>nx5085);
   ix5086 : mux21 port map ( Y=>nx5085, A0=>nx5036, A1=>nx5042, S0=>nx5038);
   ix5088 : mux21 port map ( Y=>nx5087, A0=>nx5002, A1=>nx5044, S0=>nx1893);
   ix4523 : nor02 port map ( Y=>mac_output(28), A0=>RST, A1=>nx5090);
   ix5091 : nand02 port map ( Y=>nx5090, A0=>nx2523, A1=>nx4232);
   ix4233 : xnor2 port map ( Y=>nx4232, A0=>nx1891, A1=>nx5122);
   ix4241 : xnor2 port map ( Y=>nx1891, A0=>mac_unit_tempP_28, A1=>nx5096);
   mac_unit_MR_reg_Q_28 : dffr port map ( Q=>mac_unit_tempP_28, QB=>OPEN, D
      =>nx4232, CLK=>CLK, R=>RST);
   ix5097 : xnor2 port map ( Y=>nx5096, A0=>nx5098, A1=>nx5100);
   ix5099 : mux21 port map ( Y=>nx5098, A0=>nx5055, A1=>nx5061, S0=>nx5057);
   ix5101 : xnor2 port map ( Y=>nx5100, A0=>nx5102, A1=>nx5104);
   ix5103 : nand02 port map ( Y=>nx5102, A0=>nx146, A1=>nx5520);
   ix5105 : xnor2 port map ( Y=>nx5104, A0=>nx5106, A1=>nx5108);
   ix5107 : mux21 port map ( Y=>nx5106, A0=>nx5063, A1=>nx5069, S0=>nx5065);
   ix5109 : xnor2 port map ( Y=>nx5108, A0=>nx5110, A1=>nx5112);
   ix5111 : nand02 port map ( Y=>nx5110, A0=>nx5516, A1=>nx122);
   ix5113 : xnor2 port map ( Y=>nx5112, A0=>nx5114, A1=>nx5116);
   ix5115 : mux21 port map ( Y=>nx5114, A0=>nx5071, A1=>nx5077, S0=>nx5073);
   ix5117 : xnor2 port map ( Y=>nx5116, A0=>nx5118, A1=>nx5120);
   ix5121 : mux21 port map ( Y=>nx5120, A0=>nx5079, A1=>nx5085, S0=>nx5081);
   ix5123 : mux21 port map ( Y=>nx5122, A0=>nx5053, A1=>nx5087, S0=>nx1892);
   ix4531 : nor02 port map ( Y=>mac_output(29), A0=>RST, A1=>nx5125);
   ix5126 : nand02 port map ( Y=>nx5125, A0=>nx2523, A1=>nx4250);
   ix4251 : xnor2 port map ( Y=>nx4250, A0=>nx1889, A1=>nx5149);
   ix4259 : xnor2 port map ( Y=>nx1889, A0=>mac_unit_tempP_29, A1=>nx5131);
   mac_unit_MR_reg_Q_29 : dffr port map ( Q=>mac_unit_tempP_29, QB=>OPEN, D
      =>nx4250, CLK=>CLK, R=>RST);
   ix5132 : xnor2 port map ( Y=>nx5131, A0=>nx5133, A1=>nx5135);
   ix5134 : mux21 port map ( Y=>nx5133, A0=>nx5098, A1=>nx5104, S0=>nx5100);
   ix5136 : xnor2 port map ( Y=>nx5135, A0=>nx5137, A1=>nx5139);
   ix5138 : nand02 port map ( Y=>nx5137, A0=>nx122, A1=>nx5520);
   ix5140 : xnor2 port map ( Y=>nx5139, A0=>nx5141, A1=>nx5143);
   ix5142 : mux21 port map ( Y=>nx5141, A0=>nx5106, A1=>nx5112, S0=>nx5108);
   ix5144 : xnor2 port map ( Y=>nx5143, A0=>nx5145, A1=>nx5147);
   ix5148 : mux21 port map ( Y=>nx5147, A0=>nx5114, A1=>nx5120, S0=>nx5116);
   ix5150 : mux21 port map ( Y=>nx5149, A0=>nx5096, A1=>nx5122, S0=>nx1891);
   ix4539 : nor02 port map ( Y=>mac_output(30), A0=>RST, A1=>nx5152);
   ix5153 : nand02 port map ( Y=>nx5152, A0=>nx2523, A1=>nx4268);
   ix4269 : xnor2 port map ( Y=>nx4268, A0=>nx1887, A1=>nx5168);
   ix4277 : xnor2 port map ( Y=>nx1887, A0=>mac_unit_tempP_30, A1=>nx5158);
   mac_unit_MR_reg_Q_30 : dffr port map ( Q=>mac_unit_tempP_30, QB=>OPEN, D
      =>nx4268, CLK=>CLK, R=>RST);
   ix5159 : xnor2 port map ( Y=>nx5158, A0=>nx5160, A1=>nx5162);
   ix5161 : mux21 port map ( Y=>nx5160, A0=>nx5133, A1=>nx5139, S0=>nx5135);
   ix5163 : xnor2 port map ( Y=>nx5162, A0=>nx5164, A1=>nx5166);
   ix5167 : mux21 port map ( Y=>nx5166, A0=>nx5141, A1=>nx5147, S0=>nx5143);
   ix5169 : mux21 port map ( Y=>nx5168, A0=>nx5131, A1=>nx5149, S0=>nx1889);
   ix4291 : nor02ii port map ( Y=>mac_output(31), A0=>RST, A1=>nx1885);
   ix4287 : xnor2 port map ( Y=>nx1885, A0=>nx3636, A1=>nx5177);
   ix3637 : xnor2 port map ( Y=>nx3636, A0=>mac_unit_tempP_31, A1=>nx5175);
   mac_unit_MR_reg_Q_31 : dffr port map ( Q=>mac_unit_tempP_31, QB=>OPEN, D
      =>nx1885, CLK=>CLK, R=>RST);
   ix5176 : mux21 port map ( Y=>nx5175, A0=>nx5160, A1=>nx5166, S0=>nx5162);
   ix5178 : mux21 port map ( Y=>nx5177, A0=>nx5158, A1=>nx5168, S0=>nx1887);
   test_output_reg_signature_0 : dff port map ( Q=>sig_0, QB=>OPEN, D=>
      test_output_misr_signal_31, CLK=>CLK);
   ix2416 : oai32 port map ( Y=>nx2415, A0=>nx5183, A1=>RST, A2=>nx5526, B0
      =>nx5345, B1=>nx5542);
   ix5184 : xnor2 port map ( Y=>nx5183, A0=>nx4294, A1=>
      test_output_misr_signal_30);
   ix4295 : nor02 port map ( Y=>nx4294, A0=>RST, A1=>nx2429);
   test_output_reg_misr_signal_30 : dffr port map ( Q=>
      test_output_misr_signal_30, QB=>OPEN, D=>nx2405, CLK=>CLK, R=>RST);
   ix2396 : oai32 port map ( Y=>nx2395, A0=>nx5191, A1=>RST, A2=>nx5526, B0
      =>nx5342, B1=>nx5542);
   ix2386 : oai32 port map ( Y=>nx2385, A0=>nx5195, A1=>RST, A2=>nx5526, B0
      =>nx5340, B1=>nx5542);
   ix2376 : oai32 port map ( Y=>nx2375, A0=>nx5199, A1=>RST, A2=>nx5526, B0
      =>nx5338, B1=>nx5542);
   ix2366 : oai32 port map ( Y=>nx2365, A0=>nx5203, A1=>RST, A2=>nx5526, B0
      =>nx5336, B1=>nx5542);
   ix2356 : oai32 port map ( Y=>nx2355, A0=>nx5207, A1=>RST, A2=>nx5526, B0
      =>nx5334, B1=>nx5446);
   ix2346 : oai32 port map ( Y=>nx2345, A0=>nx5211, A1=>RST, A2=>nx5526, B0
      =>nx5332, B1=>nx5446);
   ix2336 : oai32 port map ( Y=>nx2335, A0=>nx5215, A1=>RST, A2=>nx5524, B0
      =>nx5330, B1=>nx5446);
   ix2326 : oai32 port map ( Y=>nx2325, A0=>nx5219, A1=>RST, A2=>nx5524, B0
      =>nx5328, B1=>nx5446);
   ix2316 : oai32 port map ( Y=>nx2315, A0=>nx5223, A1=>RST, A2=>nx5524, B0
      =>nx5326, B1=>nx5446);
   ix2306 : oai32 port map ( Y=>nx2305, A0=>nx5227, A1=>RST, A2=>nx5524, B0
      =>nx5324, B1=>nx5446);
   ix2296 : oai32 port map ( Y=>nx2295, A0=>nx5231, A1=>RST, A2=>nx5524, B0
      =>nx5322, B1=>nx5446);
   ix2286 : oai32 port map ( Y=>nx2285, A0=>nx5235, A1=>RST, A2=>nx5524, B0
      =>nx5320, B1=>nx5446);
   ix2276 : oai32 port map ( Y=>nx2275, A0=>nx5239, A1=>RST, A2=>nx5524, B0
      =>nx5318, B1=>nx5446);
   ix2266 : oai32 port map ( Y=>nx2265, A0=>nx5243, A1=>RST, A2=>nx5524, B0
      =>nx5316, B1=>nx5446);
   ix2256 : oai32 port map ( Y=>nx2255, A0=>nx5247, A1=>RST, A2=>nx5524, B0
      =>nx5314, B1=>nx5446);
   ix5248 : xnor2 port map ( Y=>nx5247, A0=>nx4422, A1=>
      test_output_misr_signal_14);
   test_output_reg_misr_signal_14 : dffr port map ( Q=>
      test_output_misr_signal_14, QB=>OPEN, D=>nx2245, CLK=>CLK, R=>RST);
   ix2236 : oai32 port map ( Y=>nx2235, A0=>nx5254, A1=>RST, A2=>nx5524, B0
      =>nx5311, B1=>nx5446);
   ix5255 : xnor2 port map ( Y=>nx5254, A0=>nx4438, A1=>
      test_output_misr_signal_12);
   test_output_reg_misr_signal_12 : dffr port map ( Q=>
      test_output_misr_signal_12, QB=>OPEN, D=>nx2225, CLK=>CLK, R=>RST);
   ix4617 : xnor2 port map ( Y=>nx4616, A0=>nx4391, A1=>
      test_output_misr_signal_11);
   test_output_reg_misr_signal_11 : dffr port map ( Q=>
      test_output_misr_signal_11, QB=>OPEN, D=>nx2215, CLK=>CLK, R=>RST);
   ix4611 : xnor2 port map ( Y=>nx4610, A0=>nx4511, A1=>
      test_output_misr_signal_10);
   test_output_reg_misr_signal_10 : dffr port map ( Q=>
      test_output_misr_signal_10, QB=>OPEN, D=>nx2205, CLK=>CLK, R=>RST);
   ix4605 : xnor2 port map ( Y=>nx4604, A0=>nx4613, A1=>
      test_output_misr_signal_9);
   test_output_reg_misr_signal_9 : dffr port map ( Q=>
      test_output_misr_signal_9, QB=>OPEN, D=>nx2195, CLK=>CLK, R=>RST);
   ix4599 : xnor2 port map ( Y=>nx4598, A0=>nx4707, A1=>
      test_output_misr_signal_8);
   test_output_reg_misr_signal_8 : dffr port map ( Q=>
      test_output_misr_signal_8, QB=>OPEN, D=>nx2185, CLK=>CLK, R=>RST);
   ix4593 : xnor2 port map ( Y=>nx4592, A0=>nx4793, A1=>
      test_output_misr_signal_7);
   test_output_reg_misr_signal_7 : dffr port map ( Q=>
      test_output_misr_signal_7, QB=>OPEN, D=>nx2175, CLK=>CLK, R=>RST);
   ix4587 : xnor2 port map ( Y=>nx4586, A0=>nx4868, A1=>
      test_output_misr_signal_6);
   test_output_reg_misr_signal_6 : dffr port map ( Q=>
      test_output_misr_signal_6, QB=>OPEN, D=>nx2165, CLK=>CLK, R=>RST);
   ix4581 : xnor2 port map ( Y=>nx4580, A0=>nx4937, A1=>
      test_output_misr_signal_5);
   test_output_reg_misr_signal_5 : dffr port map ( Q=>
      test_output_misr_signal_5, QB=>OPEN, D=>nx2155, CLK=>CLK, R=>RST);
   ix4575 : xnor2 port map ( Y=>nx4574, A0=>nx4996, A1=>
      test_output_misr_signal_4);
   test_output_reg_misr_signal_4 : dffr port map ( Q=>
      test_output_misr_signal_4, QB=>OPEN, D=>nx2145, CLK=>CLK, R=>RST);
   ix4569 : xnor2 port map ( Y=>nx4568, A0=>nx5047, A1=>
      test_output_misr_signal_3);
   test_output_reg_misr_signal_3 : dffr port map ( Q=>
      test_output_misr_signal_3, QB=>OPEN, D=>nx2135, CLK=>CLK, R=>RST);
   ix4563 : xnor2 port map ( Y=>nx4562, A0=>nx5090, A1=>
      test_output_misr_signal_2);
   test_output_reg_misr_signal_2 : dffr port map ( Q=>
      test_output_misr_signal_2, QB=>OPEN, D=>nx2125, CLK=>CLK, R=>RST);
   ix4557 : xnor2 port map ( Y=>nx4556, A0=>nx5125, A1=>
      test_output_misr_signal_1);
   test_output_reg_misr_signal_1 : dffr port map ( Q=>
      test_output_misr_signal_1, QB=>OPEN, D=>nx2115, CLK=>CLK, R=>RST);
   ix4551 : xnor2 port map ( Y=>nx4550, A0=>nx5152, A1=>
      test_output_misr_signal_0);
   test_output_reg_misr_signal_0 : dffr port map ( Q=>
      test_output_misr_signal_0, QB=>OPEN, D=>nx2105, CLK=>CLK, R=>RST);
   ix4545 : xnor2 port map ( Y=>nx4544, A0=>nx4868, A1=>nx4542);
   test_output_reg_misr_signal_13 : dffr port map ( Q=>
      test_output_misr_signal_13, QB=>nx5311, D=>nx2235, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_15 : dffr port map ( Q=>
      test_output_misr_signal_15, QB=>nx5314, D=>nx2255, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_16 : dffr port map ( Q=>
      test_output_misr_signal_16, QB=>nx5316, D=>nx2265, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_17 : dffr port map ( Q=>
      test_output_misr_signal_17, QB=>nx5318, D=>nx2275, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_18 : dffr port map ( Q=>
      test_output_misr_signal_18, QB=>nx5320, D=>nx2285, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_19 : dffr port map ( Q=>
      test_output_misr_signal_19, QB=>nx5322, D=>nx2295, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_20 : dffr port map ( Q=>
      test_output_misr_signal_20, QB=>nx5324, D=>nx2305, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_21 : dffr port map ( Q=>
      test_output_misr_signal_21, QB=>nx5326, D=>nx2315, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_22 : dffr port map ( Q=>
      test_output_misr_signal_22, QB=>nx5328, D=>nx2325, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_23 : dffr port map ( Q=>
      test_output_misr_signal_23, QB=>nx5330, D=>nx2335, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_24 : dffr port map ( Q=>
      test_output_misr_signal_24, QB=>nx5332, D=>nx2345, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_25 : dffr port map ( Q=>
      test_output_misr_signal_25, QB=>nx5334, D=>nx2355, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_26 : dffr port map ( Q=>
      test_output_misr_signal_26, QB=>nx5336, D=>nx2365, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_27 : dffr port map ( Q=>
      test_output_misr_signal_27, QB=>nx5338, D=>nx2375, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_28 : dffr port map ( Q=>
      test_output_misr_signal_28, QB=>nx5340, D=>nx2385, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_29 : dffr port map ( Q=>
      test_output_misr_signal_29, QB=>nx5342, D=>nx2395, CLK=>CLK, R=>RST);
   test_output_reg_misr_signal_31 : dffr port map ( Q=>
      test_output_misr_signal_31, QB=>nx5345, D=>nx2415, CLK=>CLK, R=>RST);
   test_output_reg_signature_1 : dff port map ( Q=>sig_1, QB=>OPEN, D=>
      test_output_misr_signal_30, CLK=>CLK);
   test_output_reg_signature_2 : dff port map ( Q=>sig_2, QB=>OPEN, D=>
      test_output_misr_signal_29, CLK=>CLK);
   test_output_reg_signature_3 : dff port map ( Q=>sig_3, QB=>OPEN, D=>
      test_output_misr_signal_28, CLK=>CLK);
   test_output_reg_signature_4 : dff port map ( Q=>sig_4, QB=>OPEN, D=>
      test_output_misr_signal_27, CLK=>CLK);
   test_output_reg_signature_5 : dff port map ( Q=>sig_5, QB=>OPEN, D=>
      test_output_misr_signal_26, CLK=>CLK);
   test_output_reg_signature_6 : dff port map ( Q=>sig_6, QB=>OPEN, D=>
      test_output_misr_signal_25, CLK=>CLK);
   test_output_reg_signature_7 : dff port map ( Q=>sig_7, QB=>OPEN, D=>
      test_output_misr_signal_24, CLK=>CLK);
   test_output_reg_signature_8 : dff port map ( Q=>sig_8, QB=>OPEN, D=>
      test_output_misr_signal_23, CLK=>CLK);
   test_output_reg_signature_9 : dff port map ( Q=>sig_9, QB=>OPEN, D=>
      test_output_misr_signal_22, CLK=>CLK);
   test_output_reg_signature_10 : dff port map ( Q=>sig_10, QB=>OPEN, D=>
      test_output_misr_signal_21, CLK=>CLK);
   test_output_reg_signature_11 : dff port map ( Q=>sig_11, QB=>OPEN, D=>
      test_output_misr_signal_20, CLK=>CLK);
   test_output_reg_signature_12 : dff port map ( Q=>sig_12, QB=>OPEN, D=>
      test_output_misr_signal_19, CLK=>CLK);
   test_output_reg_signature_13 : dff port map ( Q=>sig_13, QB=>OPEN, D=>
      test_output_misr_signal_18, CLK=>CLK);
   test_output_reg_signature_14 : dff port map ( Q=>sig_14, QB=>OPEN, D=>
      test_output_misr_signal_17, CLK=>CLK);
   test_output_reg_signature_15 : dff port map ( Q=>sig_15, QB=>OPEN, D=>
      test_output_misr_signal_16, CLK=>CLK);
   test_output_reg_signature_16 : dff port map ( Q=>sig_16, QB=>OPEN, D=>
      test_output_misr_signal_15, CLK=>CLK);
   test_output_reg_signature_17 : dff port map ( Q=>sig_17, QB=>OPEN, D=>
      test_output_misr_signal_14, CLK=>CLK);
   test_output_reg_signature_18 : dff port map ( Q=>sig_18, QB=>OPEN, D=>
      test_output_misr_signal_13, CLK=>CLK);
   test_output_reg_signature_19 : dff port map ( Q=>sig_19, QB=>OPEN, D=>
      test_output_misr_signal_12, CLK=>CLK);
   test_output_reg_signature_20 : dff port map ( Q=>sig_20, QB=>OPEN, D=>
      test_output_misr_signal_11, CLK=>CLK);
   test_output_reg_signature_21 : dff port map ( Q=>sig_21, QB=>OPEN, D=>
      test_output_misr_signal_10, CLK=>CLK);
   test_output_reg_signature_22 : dff port map ( Q=>sig_22, QB=>OPEN, D=>
      test_output_misr_signal_9, CLK=>CLK);
   test_output_reg_signature_23 : dff port map ( Q=>sig_23, QB=>OPEN, D=>
      test_output_misr_signal_8, CLK=>CLK);
   test_output_reg_signature_24 : dff port map ( Q=>sig_24, QB=>OPEN, D=>
      test_output_misr_signal_7, CLK=>CLK);
   test_output_reg_signature_25 : dff port map ( Q=>sig_25, QB=>OPEN, D=>
      test_output_misr_signal_6, CLK=>CLK);
   test_output_reg_signature_26 : dff port map ( Q=>sig_26, QB=>OPEN, D=>
      test_output_misr_signal_5, CLK=>CLK);
   test_output_reg_signature_27 : dff port map ( Q=>sig_27, QB=>OPEN, D=>
      test_output_misr_signal_4, CLK=>CLK);
   test_output_reg_signature_28 : dff port map ( Q=>sig_28, QB=>OPEN, D=>
      test_output_misr_signal_3, CLK=>CLK);
   test_output_reg_signature_29 : dff port map ( Q=>sig_29, QB=>OPEN, D=>
      test_output_misr_signal_2, CLK=>CLK);
   test_output_reg_signature_30 : dff port map ( Q=>sig_30, QB=>OPEN, D=>
      test_output_misr_signal_1, CLK=>CLK);
   test_output_reg_signature_31 : dff port map ( Q=>sig_31, QB=>OPEN, D=>
      test_output_misr_signal_0, CLK=>CLK);
   ix4053 : inv01 port map ( Y=>nx4052, A=>nx4251);
   ix4051 : inv01 port map ( Y=>nx4050, A=>nx4257);
   ix4017 : inv01 port map ( Y=>nx4016, A=>nx3963);
   ix4015 : inv01 port map ( Y=>nx4014, A=>nx3971);
   ix3993 : inv01 port map ( Y=>nx3992, A=>nx3815);
   ix3991 : inv01 port map ( Y=>nx3990, A=>nx3823);
   ix3969 : inv01 port map ( Y=>nx3968, A=>nx3681);
   ix3967 : inv01 port map ( Y=>nx3966, A=>nx3687);
   ix3945 : inv01 port map ( Y=>nx3944, A=>nx3549);
   ix3943 : inv01 port map ( Y=>nx3942, A=>nx3557);
   ix3921 : inv01 port map ( Y=>nx3920, A=>nx3425);
   ix3919 : inv01 port map ( Y=>nx3918, A=>nx3433);
   ix3897 : inv01 port map ( Y=>nx3896, A=>nx3311);
   ix3895 : inv01 port map ( Y=>nx3894, A=>nx3319);
   ix3873 : inv01 port map ( Y=>nx3872, A=>nx3203);
   ix3871 : inv01 port map ( Y=>nx3870, A=>nx3211);
   ix3849 : inv01 port map ( Y=>nx3848, A=>nx3103);
   ix3847 : inv01 port map ( Y=>nx3846, A=>nx3111);
   ix3825 : inv01 port map ( Y=>nx3824, A=>nx3011);
   ix3823 : inv01 port map ( Y=>nx3822, A=>nx3019);
   ix3801 : inv01 port map ( Y=>nx3800, A=>nx2921);
   ix3799 : inv01 port map ( Y=>nx3798, A=>nx2929);
   ix3777 : inv01 port map ( Y=>nx3776, A=>nx2839);
   ix3775 : inv01 port map ( Y=>nx3774, A=>nx2847);
   ix3753 : inv01 port map ( Y=>nx3752, A=>nx2765);
   ix3751 : inv01 port map ( Y=>nx3750, A=>nx2773);
   ix3729 : inv01 port map ( Y=>nx3728, A=>nx2699);
   ix3727 : inv01 port map ( Y=>nx3726, A=>nx2707);
   ix3705 : inv01 port map ( Y=>nx3704, A=>nx2643);
   ix3703 : inv01 port map ( Y=>nx3702, A=>nx2651);
   ix3681 : inv01 port map ( Y=>nx3680, A=>nx2601);
   ix3679 : inv01 port map ( Y=>nx3678, A=>nx2609);
   ix3639 : inv01 port map ( Y=>nx3638, A=>nx2429);
   ix3695 : inv01 port map ( Y=>nx1933, A=>nx2603);
   ix3719 : inv01 port map ( Y=>nx1932, A=>nx2645);
   ix3743 : inv01 port map ( Y=>nx1931, A=>nx2701);
   ix3767 : inv01 port map ( Y=>nx1929, A=>nx2767);
   ix3791 : inv01 port map ( Y=>nx1927, A=>nx2841);
   ix3815 : inv01 port map ( Y=>nx1925, A=>nx2923);
   ix3839 : inv01 port map ( Y=>nx1923, A=>nx3013);
   ix3863 : inv01 port map ( Y=>nx1922, A=>nx3105);
   ix3887 : inv01 port map ( Y=>nx1921, A=>nx3205);
   ix3911 : inv01 port map ( Y=>nx1919, A=>nx3313);
   ix3935 : inv01 port map ( Y=>nx1917, A=>nx3427);
   ix3959 : inv01 port map ( Y=>nx1915, A=>nx3551);
   ix3983 : inv01 port map ( Y=>nx1913, A=>nx3683);
   ix4007 : inv01 port map ( Y=>nx1912, A=>nx3817);
   ix4025 : inv01 port map ( Y=>nx1911, A=>nx3965);
   ix4061 : inv01 port map ( Y=>nx1907, A=>nx4253);
   ix4110 : inv01 port map ( Y=>nx4109, A=>nx3574);
   ix4404 : inv01 port map ( Y=>nx4403, A=>nx3540);
   ix3956 : inv01 port map ( Y=>nx3955, A=>nx3420);
   ix4414 : inv01 port map ( Y=>nx4413, A=>nx3364);
   ix3808 : inv01 port map ( Y=>nx3807, A=>nx3198);
   ix3996 : inv01 port map ( Y=>nx3995, A=>nx3134);
   ix4128 : inv01 port map ( Y=>nx4127, A=>nx3096);
   ix4280 : inv01 port map ( Y=>nx4279, A=>nx3086);
   ix3674 : inv01 port map ( Y=>nx3673, A=>nx2976);
   ix3856 : inv01 port map ( Y=>nx3855, A=>nx2912);
   ix4138 : inv01 port map ( Y=>nx4137, A=>nx2864);
   ix4290 : inv01 port map ( Y=>nx4289, A=>nx2854);
   ix3542 : inv01 port map ( Y=>nx3541, A=>nx2754);
   ix3718 : inv01 port map ( Y=>nx3717, A=>nx2690);
   ix4148 : inv01 port map ( Y=>nx4147, A=>nx2632);
   ix4300 : inv01 port map ( Y=>nx4299, A=>nx2622);
   ix3418 : inv01 port map ( Y=>nx3417, A=>nx2532);
   ix3590 : inv01 port map ( Y=>nx3589, A=>nx2468);
   ix4158 : inv01 port map ( Y=>nx4157, A=>nx2400);
   ix4310 : inv01 port map ( Y=>nx4309, A=>nx2390);
   ix3304 : inv01 port map ( Y=>nx3303, A=>nx2310);
   ix3466 : inv01 port map ( Y=>nx3465, A=>nx2246);
   ix4168 : inv01 port map ( Y=>nx4167, A=>nx2168);
   ix4320 : inv01 port map ( Y=>nx4319, A=>nx2158);
   ix3196 : inv01 port map ( Y=>nx3195, A=>nx2088);
   ix3352 : inv01 port map ( Y=>nx3351, A=>nx2024);
   ix4178 : inv01 port map ( Y=>nx4177, A=>nx1936);
   ix4330 : inv01 port map ( Y=>nx4329, A=>nx1926);
   ix3096 : inv01 port map ( Y=>nx3095, A=>nx1866);
   ix3244 : inv01 port map ( Y=>nx3243, A=>nx1802);
   ix4188 : inv01 port map ( Y=>nx4187, A=>nx1704);
   ix4340 : inv01 port map ( Y=>nx4339, A=>nx1694);
   ix3004 : inv01 port map ( Y=>nx3003, A=>nx1644);
   ix3144 : inv01 port map ( Y=>nx3143, A=>nx1580);
   ix4198 : inv01 port map ( Y=>nx4197, A=>nx1472);
   ix4350 : inv01 port map ( Y=>nx4349, A=>nx1462);
   ix2914 : inv01 port map ( Y=>nx2913, A=>nx1422);
   ix3052 : inv01 port map ( Y=>nx3051, A=>nx1358);
   ix4206 : inv01 port map ( Y=>nx4205, A=>nx1240);
   ix4360 : inv01 port map ( Y=>nx4359, A=>nx1230);
   ix2832 : inv01 port map ( Y=>nx2831, A=>nx1200);
   ix2966 : inv01 port map ( Y=>nx2965, A=>nx1136);
   ix4216 : inv01 port map ( Y=>nx4215, A=>nx1008);
   ix4370 : inv01 port map ( Y=>nx4369, A=>nx998);
   ix2758 : inv01 port map ( Y=>nx2757, A=>nx978);
   ix2884 : inv01 port map ( Y=>nx2883, A=>nx914);
   ix4224 : inv01 port map ( Y=>nx4223, A=>nx776);
   ix4380 : inv01 port map ( Y=>nx4379, A=>nx766);
   ix2692 : inv01 port map ( Y=>nx2691, A=>nx756);
   ix2810 : inv01 port map ( Y=>nx2809, A=>nx692);
   ix4234 : inv01 port map ( Y=>nx4233, A=>nx544);
   ix2636 : inv01 port map ( Y=>nx2635, A=>nx528);
   ix4388 : inv01 port map ( Y=>nx4387, A=>nx520);
   ix2744 : inv01 port map ( Y=>nx2743, A=>nx464);
   ix2580 : inv01 port map ( Y=>nx2579, A=>nx456);
   ix2592 : inv01 port map ( Y=>nx2591, A=>nx434);
   ix2584 : inv01 port map ( Y=>nx2583, A=>nx114);
   ix4092 : inv01 port map ( Y=>nx4091, A=>nx98);
   ix2588 : inv01 port map ( Y=>nx2587, A=>nx90);
   ix5445 : inv01 port map ( Y=>nx5446, A=>nx5534);
   ix5447 : inv01 port map ( Y=>nx5448, A=>nx2587);
   ix5449 : inv01 port map ( Y=>nx5450, A=>nx2587);
   ix5455 : inv01 port map ( Y=>nx5456, A=>nx2583);
   ix5463 : inv01 port map ( Y=>nx5464, A=>nx5548);
   ix5467 : inv01 port map ( Y=>nx5468, A=>nx2635);
   ix5471 : inv01 port map ( Y=>nx5472, A=>nx2691);
   ix5475 : inv01 port map ( Y=>nx5476, A=>nx2757);
   ix5479 : inv01 port map ( Y=>nx5480, A=>nx2831);
   ix5483 : inv01 port map ( Y=>nx5484, A=>nx2913);
   ix5487 : inv01 port map ( Y=>nx5488, A=>nx3003);
   ix5491 : inv01 port map ( Y=>nx5492, A=>nx3095);
   ix5495 : inv01 port map ( Y=>nx5496, A=>nx3195);
   ix5499 : inv01 port map ( Y=>nx5500, A=>nx3303);
   ix5503 : inv01 port map ( Y=>nx5504, A=>nx3417);
   ix5507 : inv01 port map ( Y=>nx5508, A=>nx3541);
   ix5511 : inv01 port map ( Y=>nx5512, A=>nx3673);
   ix5515 : inv01 port map ( Y=>nx5516, A=>nx3807);
   ix5519 : inv01 port map ( Y=>nx5520, A=>nx3955);
   ix5523 : inv01 port map ( Y=>nx5524, A=>test_mode);
   ix5525 : inv01 port map ( Y=>nx5526, A=>test_mode);
   ix5533 : inv02 port map ( Y=>nx5534, A=>nx10);
   ix5535 : inv01 port map ( Y=>nx5536, A=>nx456);
   ix2440 : or02 port map ( Y=>nx2439, A0=>nx2587, A1=>nx5548);
   ix2096 : mux21 port map ( Y=>nx2095, A0=>test_input_lfsr_signal_15, A1=>
      test_input_lfsr_signal_14, S0=>nx5542);
   ix2086 : mux21 port map ( Y=>nx2085, A0=>test_input_lfsr_signal_14, A1=>
      test_input_lfsr_signal_13, S0=>nx5542);
   ix2076 : mux21 port map ( Y=>nx2075, A0=>test_input_lfsr_signal_13, A1=>
      test_input_lfsr_signal_12, S0=>nx5542);
   ix2066 : mux21 port map ( Y=>nx2065, A0=>test_input_lfsr_signal_12, A1=>
      test_input_lfsr_signal_11, S0=>nx5542);
   ix2056 : mux21 port map ( Y=>nx2055, A0=>test_input_lfsr_signal_11, A1=>
      test_input_lfsr_signal_10, S0=>nx5542);
   ix2046 : mux21 port map ( Y=>nx2045, A0=>test_input_lfsr_signal_10, A1=>
      test_input_lfsr_signal_9, S0=>nx5542);
   ix2036 : mux21 port map ( Y=>nx2035, A0=>test_input_lfsr_signal_9, A1=>
      test_input_lfsr_signal_8, S0=>nx5542);
   ix2026 : mux21 port map ( Y=>nx2025, A0=>test_input_lfsr_signal_8, A1=>
      test_input_lfsr_signal_7, S0=>nx5542);
   ix2016 : mux21 port map ( Y=>nx2015, A0=>test_input_lfsr_signal_7, A1=>
      test_input_lfsr_signal_6, S0=>nx5542);
   ix2006 : mux21 port map ( Y=>nx2005, A0=>test_input_lfsr_signal_6, A1=>
      test_input_lfsr_signal_5, S0=>nx5542);
   ix1996 : mux21 port map ( Y=>nx1995, A0=>test_input_lfsr_signal_5, A1=>
      test_input_lfsr_signal_4, S0=>nx5544);
   ix1986 : mux21 port map ( Y=>nx1985, A0=>test_input_lfsr_signal_4, A1=>
      test_input_lfsr_signal_3, S0=>nx5544);
   ix1976 : mux21 port map ( Y=>nx1975, A0=>test_input_lfsr_signal_3, A1=>
      test_input_lfsr_signal_2, S0=>nx5544);
   ix1966 : mux21 port map ( Y=>nx1965, A0=>test_input_lfsr_signal_2, A1=>
      test_input_lfsr_signal_1, S0=>nx5544);
   ix1956 : mux21 port map ( Y=>nx1955, A0=>test_input_lfsr_signal_1, A1=>
      test_input_lfsr_signal_0, S0=>nx5544);
   ix2522 : nor02ii port map ( Y=>nx10, A0=>RST, A1=>test_mode);
   ix2568 : or04 port map ( Y=>nx2567, A0=>nx2587, A1=>nx5548, A2=>nx2583, 
      A3=>nx2591);
   ix3665 : ao22 port map ( Y=>nx3664, A0=>nx456, A1=>nx114, B0=>nx90, B1=>
      nx434);
   ix2614 : or02 port map ( Y=>nx2613, A0=>nx5548, A1=>nx2635);
   ix2626 : or02 port map ( Y=>nx2625, A0=>nx2583, A1=>nx2591);
   ix2662 : or02 port map ( Y=>nx2661, A0=>nx5548, A1=>nx2691);
   ix2674 : or02 port map ( Y=>nx2673, A0=>nx2591, A1=>nx2635);
   ix2718 : or02 port map ( Y=>nx2717, A0=>nx5548, A1=>nx2757);
   ix2730 : or02 port map ( Y=>nx2729, A0=>nx2591, A1=>nx2691);
   ix2784 : or02 port map ( Y=>nx2783, A0=>nx5548, A1=>nx2831);
   ix2796 : or02 port map ( Y=>nx2795, A0=>nx2591, A1=>nx2757);
   ix2858 : or02 port map ( Y=>nx2857, A0=>nx5548, A1=>nx2913);
   ix2870 : or02 port map ( Y=>nx2869, A0=>nx2591, A1=>nx2831);
   ix2940 : or02 port map ( Y=>nx2939, A0=>nx5548, A1=>nx3003);
   ix2952 : or02 port map ( Y=>nx2951, A0=>nx2591, A1=>nx2913);
   ix3030 : or02 port map ( Y=>nx3029, A0=>nx5548, A1=>nx3095);
   ix3038 : or02 port map ( Y=>nx3037, A0=>nx2591, A1=>nx3003);
   ix3122 : or02 port map ( Y=>nx3121, A0=>nx5548, A1=>nx3195);
   ix3130 : or02 port map ( Y=>nx3129, A0=>nx2591, A1=>nx3095);
   ix3222 : or02 port map ( Y=>nx3221, A0=>nx5548, A1=>nx3303);
   ix3230 : or02 port map ( Y=>nx3229, A0=>nx2591, A1=>nx3195);
   ix3330 : or02 port map ( Y=>nx3329, A0=>nx5548, A1=>nx3417);
   ix3338 : or02 port map ( Y=>nx3337, A0=>nx2591, A1=>nx3303);
   ix3444 : or02 port map ( Y=>nx3443, A0=>nx5548, A1=>nx3541);
   ix3452 : or02 port map ( Y=>nx3451, A0=>nx2591, A1=>nx3417);
   ix3568 : or02 port map ( Y=>nx3567, A0=>nx5548, A1=>nx3673);
   ix3576 : or02 port map ( Y=>nx3575, A0=>nx2591, A1=>nx3541);
   ix3698 : or02 port map ( Y=>nx3697, A0=>nx2579, A1=>nx3807);
   ix3706 : or02 port map ( Y=>nx3705, A0=>nx2591, A1=>nx3673);
   ix3834 : or02 port map ( Y=>nx3833, A0=>nx2579, A1=>nx3955);
   ix3842 : or02 port map ( Y=>nx3841, A0=>nx2591, A1=>nx3807);
   ix3950 : or02 port map ( Y=>nx3949, A0=>nx2587, A1=>nx5550);
   ix3982 : or02 port map ( Y=>nx3981, A0=>nx2591, A1=>nx3955);
   ix4086 : or02 port map ( Y=>nx4085, A0=>nx2583, A1=>nx5550);
   ix4238 : or02 port map ( Y=>nx4237, A0=>nx2635, A1=>nx5550);
   ix4384 : or02 port map ( Y=>nx4383, A0=>nx2691, A1=>nx5550);
   ix4498 : or02 port map ( Y=>nx4497, A0=>nx2757, A1=>nx5550);
   ix4606 : or02 port map ( Y=>nx4605, A0=>nx2831, A1=>nx5550);
   ix4700 : or02 port map ( Y=>nx4699, A0=>nx2913, A1=>nx5550);
   ix4786 : or02 port map ( Y=>nx4785, A0=>nx3003, A1=>nx5550);
   ix4862 : or02 port map ( Y=>nx4861, A0=>nx3095, A1=>nx5550);
   ix4930 : or02 port map ( Y=>nx4929, A0=>nx3195, A1=>nx5550);
   ix4990 : or02 port map ( Y=>nx4989, A0=>nx3303, A1=>nx5550);
   ix5041 : or02 port map ( Y=>nx5040, A0=>nx3417, A1=>nx5550);
   ix5084 : or02 port map ( Y=>nx5083, A0=>nx3541, A1=>nx5550);
   ix5119 : or02 port map ( Y=>nx5118, A0=>nx3673, A1=>nx5550);
   ix5146 : or02 port map ( Y=>nx5145, A0=>nx3807, A1=>nx4091);
   ix5165 : or02 port map ( Y=>nx5164, A0=>nx3955, A1=>nx4091);
   ix4743 : and02 port map ( Y=>signature(0), A0=>test_mode, A1=>sig_0);
   ix2406 : mux21 port map ( Y=>nx2405, A0=>test_output_misr_signal_30, A1=>
      nx4724, S0=>nx5544);
   ix4725 : xor2 port map ( Y=>nx4724, A0=>nx2555, A1=>nx5342);
   ix5192 : xor2 port map ( Y=>nx5191, A0=>nx4310, A1=>nx5340);
   ix5196 : xor2 port map ( Y=>nx5195, A0=>nx4318, A1=>nx5338);
   ix5200 : xor2 port map ( Y=>nx5199, A0=>nx4326, A1=>nx5336);
   ix5204 : xor2 port map ( Y=>nx5203, A0=>nx4334, A1=>nx5334);
   ix5208 : xor2 port map ( Y=>nx5207, A0=>nx4342, A1=>nx5332);
   ix5212 : xor2 port map ( Y=>nx5211, A0=>nx4350, A1=>nx5330);
   ix5216 : xor2 port map ( Y=>nx5215, A0=>nx4358, A1=>nx5328);
   ix5220 : xor2 port map ( Y=>nx5219, A0=>nx4366, A1=>nx5326);
   ix5224 : xor2 port map ( Y=>nx5223, A0=>nx4374, A1=>nx5324);
   ix5228 : xor2 port map ( Y=>nx5227, A0=>nx4382, A1=>nx5322);
   ix5232 : xor2 port map ( Y=>nx5231, A0=>nx4390, A1=>nx5320);
   ix5236 : xor2 port map ( Y=>nx5235, A0=>nx4398, A1=>nx5318);
   ix5240 : xor2 port map ( Y=>nx5239, A0=>nx4406, A1=>nx5316);
   ix5244 : xor2 port map ( Y=>nx5243, A0=>nx4414, A1=>nx5314);
   ix2246 : mux21 port map ( Y=>nx2245, A0=>test_output_misr_signal_14, A1=>
      nx4628, S0=>nx5544);
   ix4629 : xor2 port map ( Y=>nx4628, A0=>nx4095, A1=>nx5311);
   ix2226 : mux21 port map ( Y=>nx2225, A0=>test_output_misr_signal_12, A1=>
      nx4616, S0=>nx5544);
   ix2216 : mux21 port map ( Y=>nx2215, A0=>test_output_misr_signal_11, A1=>
      nx4610, S0=>nx5544);
   ix2206 : mux21 port map ( Y=>nx2205, A0=>test_output_misr_signal_10, A1=>
      nx4604, S0=>nx5544);
   ix2196 : mux21 port map ( Y=>nx2195, A0=>test_output_misr_signal_9, A1=>
      nx4598, S0=>nx5544);
   ix2186 : mux21 port map ( Y=>nx2185, A0=>test_output_misr_signal_8, A1=>
      nx4592, S0=>nx5544);
   ix2176 : mux21 port map ( Y=>nx2175, A0=>test_output_misr_signal_7, A1=>
      nx4586, S0=>nx5544);
   ix2166 : mux21 port map ( Y=>nx2165, A0=>test_output_misr_signal_6, A1=>
      nx4580, S0=>nx5544);
   ix2156 : mux21 port map ( Y=>nx2155, A0=>test_output_misr_signal_5, A1=>
      nx4574, S0=>nx5544);
   ix2146 : mux21 port map ( Y=>nx2145, A0=>test_output_misr_signal_4, A1=>
      nx4568, S0=>nx5546);
   ix2136 : mux21 port map ( Y=>nx2135, A0=>test_output_misr_signal_3, A1=>
      nx4562, S0=>nx5546);
   ix2126 : mux21 port map ( Y=>nx2125, A0=>test_output_misr_signal_2, A1=>
      nx4556, S0=>nx5546);
   ix2116 : mux21 port map ( Y=>nx2115, A0=>test_output_misr_signal_1, A1=>
      nx4550, S0=>nx5546);
   ix2106 : mux21 port map ( Y=>nx2105, A0=>test_output_misr_signal_0, A1=>
      nx4544, S0=>nx5546);
   ix4543 : xor2 port map ( Y=>nx4542, A0=>nx5334, A1=>nx5296);
   ix5297 : xnor2 port map ( Y=>nx5296, A0=>nx5345, A1=>nx5342);
   ix4751 : and02 port map ( Y=>signature(1), A0=>test_mode, A1=>sig_1);
   ix4759 : and02 port map ( Y=>signature(2), A0=>test_mode, A1=>sig_2);
   ix4767 : and02 port map ( Y=>signature(3), A0=>test_mode, A1=>sig_3);
   ix4775 : and02 port map ( Y=>signature(4), A0=>test_mode, A1=>sig_4);
   ix4783 : and02 port map ( Y=>signature(5), A0=>test_mode, A1=>sig_5);
   ix4791 : and02 port map ( Y=>signature(6), A0=>test_mode, A1=>sig_6);
   ix4799 : and02 port map ( Y=>signature(7), A0=>test_mode, A1=>sig_7);
   ix4807 : and02 port map ( Y=>signature(8), A0=>test_mode, A1=>sig_8);
   ix4815 : and02 port map ( Y=>signature(9), A0=>test_mode, A1=>sig_9);
   ix4823 : and02 port map ( Y=>signature(10), A0=>test_mode, A1=>sig_10);
   ix4831 : and02 port map ( Y=>signature(11), A0=>test_mode, A1=>sig_11);
   ix4839 : and02 port map ( Y=>signature(12), A0=>test_mode, A1=>sig_12);
   ix4847 : and02 port map ( Y=>signature(13), A0=>test_mode, A1=>sig_13);
   ix4855 : and02 port map ( Y=>signature(14), A0=>test_mode, A1=>sig_14);
   ix4863 : and02 port map ( Y=>signature(15), A0=>test_mode, A1=>sig_15);
   ix4871 : and02 port map ( Y=>signature(16), A0=>test_mode, A1=>sig_16);
   ix4879 : and02 port map ( Y=>signature(17), A0=>test_mode, A1=>sig_17);
   ix4887 : and02 port map ( Y=>signature(18), A0=>test_mode, A1=>sig_18);
   ix4895 : and02 port map ( Y=>signature(19), A0=>test_mode, A1=>sig_19);
   ix4903 : and02 port map ( Y=>signature(20), A0=>test_mode, A1=>sig_20);
   ix4911 : and02 port map ( Y=>signature(21), A0=>test_mode, A1=>sig_21);
   ix4919 : and02 port map ( Y=>signature(22), A0=>test_mode, A1=>sig_22);
   ix4927 : and02 port map ( Y=>signature(23), A0=>test_mode, A1=>sig_23);
   ix4935 : and02 port map ( Y=>signature(24), A0=>test_mode, A1=>sig_24);
   ix4943 : and02 port map ( Y=>signature(25), A0=>test_mode, A1=>sig_25);
   ix4951 : and02 port map ( Y=>signature(26), A0=>test_mode, A1=>sig_26);
   ix4959 : and02 port map ( Y=>signature(27), A0=>test_mode, A1=>sig_27);
   ix4967 : and02 port map ( Y=>signature(28), A0=>test_mode, A1=>sig_28);
   ix4975 : and02 port map ( Y=>signature(29), A0=>test_mode, A1=>sig_29);
   ix4983 : and02 port map ( Y=>signature(30), A0=>test_mode, A1=>sig_30);
   ix4991 : and02 port map ( Y=>signature(31), A0=>test_mode, A1=>sig_31);
   ix5541 : inv02 port map ( Y=>nx5542, A=>nx5534);
   ix5543 : inv02 port map ( Y=>nx5544, A=>nx5534);
   ix5545 : inv02 port map ( Y=>nx5546, A=>nx5534);
   ix5547 : inv01 port map ( Y=>nx5548, A=>nx456);
   ix5549 : inv01 port map ( Y=>nx5550, A=>nx98);
end behavioral ;

