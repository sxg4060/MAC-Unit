//
// Verilog description for cell BIST, 
// Fri Dec  6 15:00:32 2019
//
// LeonardoSpectrum Level 3, 2008b.3 
//


module BIST ( B, C, Cin, CLK, RST, test_mode, signature, mac_output ) ;

    input [15:0]B ;
    input [15:0]C ;
    input Cin ;
    input CLK ;
    input RST ;
    input test_mode ;
    output [31:0]signature ;
    output [31:0]mac_output ;

    wire mac_unit_tempP_31, nx1885, lfsr_C_15, test_input_lfsr_signal_15, nx10, 
         test_input_lfsr_signal_14, test_input_lfsr_signal_13, 
         test_input_lfsr_signal_12, test_input_lfsr_signal_11, 
         test_input_lfsr_signal_10, test_input_lfsr_signal_9, 
         test_input_lfsr_signal_8, test_input_lfsr_signal_7, 
         test_input_lfsr_signal_6, test_input_lfsr_signal_5, 
         test_input_lfsr_signal_4, test_input_lfsr_signal_3, 
         test_input_lfsr_signal_2, test_input_lfsr_signal_1, 
         test_input_lfsr_signal_0, nx14, nx90, nx98, lfsr_C_14, nx114, nx122, 
         lfsr_C_13, nx146, lfsr_C_12, nx170, lfsr_C_11, nx194, lfsr_C_10, nx218, 
         lfsr_C_9, nx242, lfsr_C_8, nx266, lfsr_C_7, nx290, lfsr_C_6, nx314, 
         lfsr_C_5, nx338, lfsr_C_4, nx362, lfsr_C_3, nx386, lfsr_C_2, nx410, 
         lfsr_C_1, nx434, lfsr_B_15, nx456, nx464, nx520, nx528, nx532, nx544, 
         nx548, nx674, nx678, nx688, nx692, nx756, nx766, nx770, nx776, nx780, 
         nx896, nx900, nx910, nx914, nx978, nx998, nx1002, nx1008, nx1012, 
         nx1118, nx1122, nx1132, nx1136, nx1200, nx1230, nx1234, nx1240, nx1244, 
         nx1340, nx1344, nx1354, nx1358, nx1422, nx1462, nx1466, nx1472, nx1476, 
         nx1562, nx1566, nx1576, nx1580, nx1644, nx1694, nx1698, nx1704, nx1708, 
         nx1784, nx1788, nx1798, nx1802, nx1866, nx1926, nx1930, nx1936, nx1940, 
         nx2006, nx2010, nx2020, nx2024, nx2088, nx2158, nx2162, nx2168, nx2172, 
         nx2228, nx2232, nx2242, nx2246, nx2310, nx2390, nx2394, nx2400, nx2404, 
         nx2450, nx2454, nx2464, nx2468, nx2532, nx2622, nx2626, nx2632, nx2636, 
         nx2672, nx2676, nx2686, nx2690, nx2754, nx2854, nx2858, nx2864, nx2868, 
         nx2894, nx2898, nx2908, nx2912, nx2976, nx3086, nx3090, nx3096, nx3100, 
         nx3116, nx3120, nx3130, nx3134, nx3198, nx3318, nx3322, nx3328, nx3332, 
         nx3338, nx3342, nx3352, nx3356, nx3360, nx3364, nx3420, nx3540, nx3544, 
         nx3574, nx3636, mac_unit_tempP_30, nx1887, mac_unit_tempP_29, nx1889, 
         mac_unit_tempP_28, nx1891, mac_unit_tempP_27, nx1892, mac_unit_tempP_26, 
         nx1893, mac_unit_tempP_25, nx1895, mac_unit_tempP_24, nx1897, 
         mac_unit_tempP_23, nx1899, mac_unit_tempP_22, nx1901, mac_unit_tempP_21, 
         nx1902, mac_unit_tempP_20, nx1903, mac_unit_tempP_19, nx1905, 
         mac_unit_tempP_18, nx1907, mac_unit_tempP_17, nx1909, mac_unit_tempP_16, 
         nx1911, mac_unit_tempP_15, nx1912, mac_unit_tempP_14, nx1913, 
         mac_unit_tempP_13, nx1915, mac_unit_tempP_12, nx1917, mac_unit_tempP_11, 
         nx1919, mac_unit_tempP_10, nx1921, mac_unit_tempP_9, nx1922, 
         mac_unit_tempP_8, nx1923, mac_unit_tempP_7, nx1925, mac_unit_tempP_6, 
         nx1927, mac_unit_tempP_5, nx1929, mac_unit_tempP_4, nx1931, 
         mac_unit_tempP_3, nx1932, mac_unit_tempP_2, nx1933, mac_unit_tempP_1, 
         nx1935, mac_unit_tempP_0, nx1937, nx3638, nx3654, nx3664, nx3678, 
         nx3680, nx3692, nx3702, nx3704, nx3716, nx3726, nx3728, nx3740, nx3750, 
         nx3752, nx3764, nx3774, nx3776, nx3788, nx3798, nx3800, nx3812, nx3822, 
         nx3824, nx3836, nx3846, nx3848, nx3860, nx3870, nx3872, nx3884, nx3894, 
         nx3896, nx3908, nx3918, nx3920, nx3932, nx3942, nx3944, nx3956, nx3966, 
         nx3968, nx3980, nx3990, nx3992, nx4004, nx4014, nx4016, nx4022, nx4034, 
         nx4050, nx4052, nx4058, nx4070, nx4088, nx4106, nx4124, nx4142, nx4160, 
         nx4178, nx4196, nx4214, nx4232, nx4250, nx4268, nx4294, nx4310, nx4318, 
         nx4326, nx4334, nx4342, nx4350, nx4358, nx4366, nx4374, nx4382, nx4390, 
         nx4398, nx4406, nx4414, nx4422, nx4438, sig_0, 
         test_output_misr_signal_31, test_output_misr_signal_30, 
         test_output_misr_signal_29, test_output_misr_signal_28, 
         test_output_misr_signal_27, test_output_misr_signal_26, 
         test_output_misr_signal_25, test_output_misr_signal_24, 
         test_output_misr_signal_23, test_output_misr_signal_22, 
         test_output_misr_signal_21, test_output_misr_signal_20, 
         test_output_misr_signal_19, test_output_misr_signal_18, 
         test_output_misr_signal_17, test_output_misr_signal_16, 
         test_output_misr_signal_15, test_output_misr_signal_14, 
         test_output_misr_signal_13, test_output_misr_signal_12, 
         test_output_misr_signal_11, test_output_misr_signal_10, 
         test_output_misr_signal_9, test_output_misr_signal_8, 
         test_output_misr_signal_7, test_output_misr_signal_6, 
         test_output_misr_signal_5, test_output_misr_signal_4, 
         test_output_misr_signal_3, test_output_misr_signal_2, 
         test_output_misr_signal_1, test_output_misr_signal_0, nx4542, nx4544, 
         nx4550, nx4556, nx4562, nx4568, nx4574, nx4580, nx4586, nx4592, nx4598, 
         nx4604, nx4610, nx4616, nx4628, nx4724, sig_1, sig_2, sig_3, sig_4, 
         sig_5, sig_6, sig_7, sig_8, sig_9, sig_10, sig_11, sig_12, sig_13, 
         sig_14, sig_15, sig_16, sig_17, sig_18, sig_19, sig_20, sig_21, sig_22, 
         sig_23, sig_24, sig_25, sig_26, sig_27, sig_28, sig_29, sig_30, sig_31, 
         nx1945, nx1955, nx1965, nx1975, nx1985, nx1995, nx2005, nx2015, nx2025, 
         nx2035, nx2045, nx2055, nx2065, nx2075, nx2085, nx2095, nx2105, nx2115, 
         nx2125, nx2135, nx2145, nx2155, nx2165, nx2175, nx2185, nx2195, nx2205, 
         nx2215, nx2225, nx2235, nx2245, nx2255, nx2265, nx2275, nx2285, nx2295, 
         nx2305, nx2315, nx2325, nx2335, nx2345, nx2355, nx2365, nx2375, nx2385, 
         nx2395, nx2405, nx2415, nx2429, nx2439, nx2509, nx2513, nx2517, nx2523, 
         nx2555, nx2565, nx2567, nx2579, nx2583, nx2587, nx2591, nx2595, nx2601, 
         nx2603, nx2609, nx2613, nx2621, nx2623, nx2625, nx2627, nx2635, nx2643, 
         nx2645, nx2651, nx2661, nx2668, nx2673, nx2679, nx2681, nx2683, nx2691, 
         nx2699, nx2701, nx2707, nx2717, nx2725, nx2729, nx2735, nx2737, nx2739, 
         nx2741, nx2743, nx2745, nx2747, nx2749, nx2757, nx2765, nx2767, nx2773, 
         nx2783, nx2790, nx2795, nx2801, nx2803, nx2805, nx2807, nx2809, nx2811, 
         nx2813, nx2815, nx2817, nx2819, nx2821, nx2823, nx2831, nx2839, nx2841, 
         nx2847, nx2857, nx2865, nx2869, nx2875, nx2877, nx2879, nx2881, nx2883, 
         nx2885, nx2887, nx2889, nx2891, nx2893, nx2895, nx2897, nx2899, nx2901, 
         nx2903, nx2905, nx2913, nx2921, nx2923, nx2929, nx2939, nx2947, nx2951, 
         nx2957, nx2959, nx2961, nx2963, nx2965, nx2967, nx2969, nx2971, nx2973, 
         nx2975, nx2977, nx2979, nx2981, nx2983, nx2985, nx2987, nx2989, nx2991, 
         nx2993, nx2995, nx3003, nx3011, nx3013, nx3019, nx3029, nx3033, nx3037, 
         nx3043, nx3045, nx3047, nx3049, nx3051, nx3053, nx3055, nx3057, nx3059, 
         nx3061, nx3063, nx3065, nx3067, nx3069, nx3071, nx3073, nx3075, nx3077, 
         nx3079, nx3081, nx3083, nx3085, nx3087, nx3089, nx3095, nx3103, nx3105, 
         nx3111, nx3121, nx3125, nx3129, nx3135, nx3137, nx3139, nx3141, nx3143, 
         nx3145, nx3147, nx3149, nx3151, nx3153, nx3155, nx3157, nx3159, nx3161, 
         nx3163, nx3165, nx3167, nx3169, nx3171, nx3173, nx3175, nx3177, nx3179, 
         nx3181, nx3183, nx3185, nx3187, nx3189, nx3195, nx3203, nx3205, nx3211, 
         nx3221, nx3225, nx3229, nx3235, nx3237, nx3239, nx3241, nx3243, nx3245, 
         nx3247, nx3249, nx3251, nx3253, nx3255, nx3257, nx3259, nx3261, nx3263, 
         nx3265, nx3267, nx3269, nx3271, nx3273, nx3275, nx3277, nx3279, nx3281, 
         nx3283, nx3285, nx3287, nx3289, nx3291, nx3293, nx3295, nx3297, nx3303, 
         nx3311, nx3313, nx3319, nx3329, nx3333, nx3337, nx3343, nx3345, nx3347, 
         nx3349, nx3351, nx3353, nx3355, nx3357, nx3359, nx3361, nx3363, nx3365, 
         nx3367, nx3369, nx3371, nx3373, nx3375, nx3377, nx3379, nx3381, nx3383, 
         nx3385, nx3387, nx3389, nx3391, nx3393, nx3395, nx3397, nx3399, nx3401, 
         nx3403, nx3405, nx3407, nx3409, nx3411, nx3413, nx3417, nx3425, nx3427, 
         nx3433, nx3443, nx3447, nx3451, nx3457, nx3459, nx3461, nx3463, nx3465, 
         nx3467, nx3469, nx3471, nx3473, nx3475, nx3477, nx3479, nx3481, nx3483, 
         nx3485, nx3487, nx3489, nx3491, nx3493, nx3495, nx3497, nx3499, nx3501, 
         nx3503, nx3505, nx3507, nx3509, nx3511, nx3513, nx3515, nx3517, nx3519, 
         nx3521, nx3523, nx3525, nx3527, nx3529, nx3531, nx3533, nx3535, nx3541, 
         nx3549, nx3551, nx3557, nx3567, nx3571, nx3575, nx3581, nx3583, nx3585, 
         nx3587, nx3589, nx3591, nx3593, nx3595, nx3597, nx3599, nx3601, nx3603, 
         nx3605, nx3607, nx3609, nx3611, nx3613, nx3615, nx3617, nx3619, nx3621, 
         nx3623, nx3625, nx3627, nx3629, nx3631, nx3633, nx3635, nx3637, nx3639, 
         nx3641, nx3643, nx3645, nx3647, nx3649, nx3651, nx3653, nx3655, nx3657, 
         nx3659, nx3661, nx3663, nx3665, nx3667, nx3673, nx3681, nx3683, nx3687, 
         nx3697, nx3701, nx3705, nx3709, nx3711, nx3713, nx3715, nx3717, nx3719, 
         nx3721, nx3723, nx3725, nx3727, nx3729, nx3731, nx3733, nx3735, nx3737, 
         nx3739, nx3741, nx3743, nx3745, nx3747, nx3749, nx3751, nx3753, nx3755, 
         nx3757, nx3759, nx3761, nx3763, nx3765, nx3767, nx3769, nx3771, nx3773, 
         nx3775, nx3777, nx3779, nx3781, nx3783, nx3785, nx3787, nx3789, nx3791, 
         nx3793, nx3795, nx3797, nx3799, nx3801, nx3803, nx3807, nx3815, nx3817, 
         nx3823, nx3833, nx3837, nx3841, nx3847, nx3849, nx3851, nx3853, nx3855, 
         nx3857, nx3859, nx3861, nx3863, nx3865, nx3867, nx3869, nx3871, nx3873, 
         nx3875, nx3877, nx3879, nx3881, nx3883, nx3885, nx3887, nx3889, nx3891, 
         nx3893, nx3895, nx3897, nx3899, nx3901, nx3903, nx3905, nx3907, nx3909, 
         nx3911, nx3913, nx3915, nx3917, nx3919, nx3921, nx3923, nx3925, nx3927, 
         nx3929, nx3931, nx3933, nx3935, nx3937, nx3939, nx3941, nx3943, nx3945, 
         nx3947, nx3949, nx3955, nx3963, nx3965, nx3971, nx3979, nx3981, nx3983, 
         nx3989, nx3993, nx3995, nx3999, nx4003, nx4007, nx4011, nx4015, nx4019, 
         nx4023, nx4027, nx4031, nx4035, nx4038, nx4041, nx4045, nx4049, nx4053, 
         nx4056, nx4059, nx4063, nx4067, nx4071, nx4074, nx4077, nx4081, nx4085, 
         nx4087, nx4091, nx4095, nx4105, nx4107, nx4109, nx4111, nx4113, nx4115, 
         nx4121, nx4125, nx4127, nx4131, nx4135, nx4137, nx4141, nx4145, nx4147, 
         nx4151, nx4155, nx4157, nx4161, nx4164, nx4167, nx4171, nx4175, nx4177, 
         nx4181, nx4185, nx4187, nx4191, nx4195, nx4197, nx4200, nx4203, nx4205, 
         nx4209, nx4213, nx4215, nx4218, nx4221, nx4223, nx4227, nx4231, nx4233, 
         nx4237, nx4239, nx4251, nx4253, nx4257, nx4261, nx4265, nx4271, nx4273, 
         nx4275, nx4277, nx4279, nx4281, nx4283, nx4285, nx4287, nx4289, nx4291, 
         nx4293, nx4295, nx4297, nx4299, nx4301, nx4303, nx4305, nx4307, nx4309, 
         nx4311, nx4313, nx4315, nx4317, nx4319, nx4321, nx4323, nx4325, nx4327, 
         nx4329, nx4331, nx4333, nx4335, nx4337, nx4339, nx4341, nx4343, nx4345, 
         nx4347, nx4349, nx4351, nx4353, nx4355, nx4357, nx4359, nx4361, nx4363, 
         nx4365, nx4367, nx4369, nx4371, nx4373, nx4375, nx4377, nx4379, nx4381, 
         nx4383, nx4385, nx4387, nx4391, nx4399, nx4401, nx4403, nx4405, nx4407, 
         nx4409, nx4411, nx4413, nx4415, nx4417, nx4419, nx4421, nx4423, nx4425, 
         nx4427, nx4429, nx4431, nx4433, nx4435, nx4437, nx4439, nx4441, nx4443, 
         nx4445, nx4447, nx4449, nx4451, nx4453, nx4455, nx4457, nx4459, nx4461, 
         nx4463, nx4465, nx4467, nx4469, nx4471, nx4473, nx4475, nx4477, nx4479, 
         nx4481, nx4483, nx4485, nx4487, nx4489, nx4491, nx4493, nx4495, nx4497, 
         nx4499, nx4501, nx4511, nx4519, nx4521, nx4523, nx4525, nx4527, nx4529, 
         nx4531, nx4533, nx4535, nx4537, nx4539, nx4541, nx4543, nx4545, nx4547, 
         nx4549, nx4551, nx4553, nx4555, nx4557, nx4559, nx4561, nx4563, nx4565, 
         nx4567, nx4569, nx4571, nx4573, nx4575, nx4577, nx4579, nx4581, nx4583, 
         nx4585, nx4587, nx4589, nx4591, nx4593, nx4595, nx4597, nx4599, nx4601, 
         nx4603, nx4605, nx4607, nx4609, nx4613, nx4620, nx4623, nx4625, nx4627, 
         nx4629, nx4631, nx4633, nx4635, nx4637, nx4639, nx4641, nx4643, nx4645, 
         nx4647, nx4649, nx4651, nx4653, nx4655, nx4657, nx4659, nx4661, nx4663, 
         nx4665, nx4667, nx4669, nx4671, nx4673, nx4675, nx4677, nx4679, nx4681, 
         nx4683, nx4685, nx4687, nx4689, nx4691, nx4693, nx4695, nx4697, nx4699, 
         nx4701, nx4703, nx4707, nx4714, nx4716, nx4719, nx4721, nx4723, nx4725, 
         nx4727, nx4729, nx4731, nx4733, nx4735, nx4737, nx4739, nx4741, nx4743, 
         nx4745, nx4747, nx4749, nx4751, nx4753, nx4755, nx4757, nx4759, nx4761, 
         nx4763, nx4765, nx4767, nx4769, nx4771, nx4773, nx4775, nx4777, nx4779, 
         nx4781, nx4783, nx4785, nx4787, nx4789, nx4793, nx4799, nx4801, nx4803, 
         nx4805, nx4807, nx4809, nx4811, nx4813, nx4815, nx4817, nx4819, nx4821, 
         nx4823, nx4825, nx4827, nx4829, nx4831, nx4833, nx4835, nx4837, nx4839, 
         nx4841, nx4843, nx4845, nx4847, nx4849, nx4851, nx4853, nx4855, nx4857, 
         nx4859, nx4861, nx4863, nx4865, nx4868, nx4875, nx4877, nx4879, nx4881, 
         nx4883, nx4885, nx4887, nx4889, nx4891, nx4893, nx4895, nx4897, nx4899, 
         nx4901, nx4903, nx4905, nx4907, nx4909, nx4911, nx4913, nx4915, nx4917, 
         nx4919, nx4921, nx4923, nx4925, nx4927, nx4929, nx4931, nx4933, nx4937, 
         nx4943, nx4945, nx4947, nx4949, nx4951, nx4953, nx4955, nx4957, nx4959, 
         nx4961, nx4963, nx4965, nx4967, nx4969, nx4971, nx4973, nx4975, nx4977, 
         nx4979, nx4981, nx4983, nx4985, nx4987, nx4989, nx4991, nx4993, nx4996, 
         nx5002, nx5004, nx5006, nx5008, nx5010, nx5012, nx5014, nx5016, nx5018, 
         nx5020, nx5022, nx5024, nx5026, nx5028, nx5030, nx5032, nx5034, nx5036, 
         nx5038, nx5040, nx5042, nx5044, nx5047, nx5053, nx5055, nx5057, nx5059, 
         nx5061, nx5063, nx5065, nx5067, nx5069, nx5071, nx5073, nx5075, nx5077, 
         nx5079, nx5081, nx5083, nx5085, nx5087, nx5090, nx5096, nx5098, nx5100, 
         nx5102, nx5104, nx5106, nx5108, nx5110, nx5112, nx5114, nx5116, nx5118, 
         nx5120, nx5122, nx5125, nx5131, nx5133, nx5135, nx5137, nx5139, nx5141, 
         nx5143, nx5145, nx5147, nx5149, nx5152, nx5158, nx5160, nx5162, nx5164, 
         nx5166, nx5168, nx5175, nx5177, nx5183, nx5191, nx5195, nx5199, nx5203, 
         nx5207, nx5211, nx5215, nx5219, nx5223, nx5227, nx5231, nx5235, nx5239, 
         nx5243, nx5247, nx5254, nx5296, nx5311, nx5314, nx5316, nx5318, nx5320, 
         nx5322, nx5324, nx5326, nx5328, nx5330, nx5332, nx5334, nx5336, nx5338, 
         nx5340, nx5342, nx5345, nx5446, nx5448, nx5450, nx5456, nx5464, nx5468, 
         nx5472, nx5476, nx5480, nx5484, nx5488, nx5492, nx5496, nx5500, nx5504, 
         nx5508, nx5512, nx5516, nx5520, nx5524, nx5526, nx5534, nx5536, nx5542, 
         nx5544, nx5546, nx5548, nx5550;
    wire [109:0] \$dummy ;




    nor02 ix4299 (.Y (mac_output[0]), .A0 (RST), .A1 (nx2429)) ;
    xnor2 ix2430 (.Y (nx2429), .A0 (Cin), .A1 (nx1937)) ;
    xnor2 ix3645 (.Y (nx1937), .A0 (mac_unit_tempP_0), .A1 (nx2439)) ;
    dffr mac_unit_MR_reg_Q_0 (.Q (mac_unit_tempP_0), .QB (\$dummy [0]), .D (
         nx3638), .CLK (CLK), .R (RST)) ;
    mux21 ix91 (.Y (nx90), .A0 (B[0]), .A1 (lfsr_C_15), .S0 (test_mode)) ;
    dff test_input_reg_BP2_15 (.Q (lfsr_C_15), .QB (\$dummy [1]), .D (
        test_input_lfsr_signal_15), .CLK (CLK)) ;
    dffs test_input_reg_lfsr_signal_15 (.Q (test_input_lfsr_signal_15), .QB (
         \$dummy [2]), .D (nx2095), .CLK (CLK), .S (RST)) ;
    dffr test_input_reg_lfsr_signal_14 (.Q (test_input_lfsr_signal_14), .QB (
         \$dummy [3]), .D (nx2085), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_13 (.Q (test_input_lfsr_signal_13), .QB (
         \$dummy [4]), .D (nx2075), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_12 (.Q (test_input_lfsr_signal_12), .QB (
         \$dummy [5]), .D (nx2065), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_11 (.Q (test_input_lfsr_signal_11), .QB (
         \$dummy [6]), .D (nx2055), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_10 (.Q (test_input_lfsr_signal_10), .QB (
         \$dummy [7]), .D (nx2045), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_9 (.Q (test_input_lfsr_signal_9), .QB (
         \$dummy [8]), .D (nx2035), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_8 (.Q (test_input_lfsr_signal_8), .QB (
         \$dummy [9]), .D (nx2025), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_7 (.Q (test_input_lfsr_signal_7), .QB (
         \$dummy [10]), .D (nx2015), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_6 (.Q (test_input_lfsr_signal_6), .QB (
         \$dummy [11]), .D (nx2005), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_5 (.Q (test_input_lfsr_signal_5), .QB (
         \$dummy [12]), .D (nx1995), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_4 (.Q (test_input_lfsr_signal_4), .QB (
         \$dummy [13]), .D (nx1985), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_3 (.Q (test_input_lfsr_signal_3), .QB (
         \$dummy [14]), .D (nx1975), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_2 (.Q (test_input_lfsr_signal_2), .QB (
         \$dummy [15]), .D (nx1965), .CLK (CLK), .R (RST)) ;
    dffr test_input_reg_lfsr_signal_1 (.Q (test_input_lfsr_signal_1), .QB (
         \$dummy [16]), .D (nx1955), .CLK (CLK), .R (RST)) ;
    oai32 ix1946 (.Y (nx1945), .A0 (nx2509), .A1 (RST), .A2 (nx5524), .B0 (
          nx2517), .B1 (nx5446)) ;
    xnor2 ix2510 (.Y (nx2509), .A0 (test_input_lfsr_signal_10), .A1 (nx14)) ;
    xnor2 ix15 (.Y (nx14), .A0 (test_input_lfsr_signal_12), .A1 (nx2513)) ;
    xnor2 ix2514 (.Y (nx2513), .A0 (test_input_lfsr_signal_15), .A1 (
          test_input_lfsr_signal_13)) ;
    dffr test_input_reg_lfsr_signal_0 (.Q (test_input_lfsr_signal_0), .QB (
         nx2517), .D (nx1945), .CLK (CLK), .R (RST)) ;
    inv01 ix2524 (.Y (nx2523), .A (RST)) ;
    mux21 ix457 (.Y (nx456), .A0 (C[0]), .A1 (lfsr_B_15), .S0 (test_mode)) ;
    dff test_input_reg_BP1_15 (.Q (lfsr_B_15), .QB (\$dummy [17]), .D (
        test_input_lfsr_signal_0), .CLK (CLK)) ;
    nor02 ix4307 (.Y (mac_output[1]), .A0 (RST), .A1 (nx2555)) ;
    nand02 ix2556 (.Y (nx2555), .A0 (nx2523), .A1 (nx3654)) ;
    xnor2 ix3655 (.Y (nx3654), .A0 (nx1935), .A1 (nx2595)) ;
    xnor2 ix3671 (.Y (nx1935), .A0 (mac_unit_tempP_1), .A1 (nx2565)) ;
    dffr mac_unit_MR_reg_Q_1 (.Q (mac_unit_tempP_1), .QB (\$dummy [18]), .D (
         nx3654), .CLK (CLK), .R (RST)) ;
    nand02 ix2566 (.Y (nx2565), .A0 (nx2567), .A1 (nx3664)) ;
    mux21 ix115 (.Y (nx114), .A0 (B[1]), .A1 (lfsr_C_14), .S0 (test_mode)) ;
    dff test_input_reg_BP2_14 (.Q (lfsr_C_14), .QB (\$dummy [19]), .D (
        test_input_lfsr_signal_14), .CLK (CLK)) ;
    mux21 ix435 (.Y (nx434), .A0 (C[1]), .A1 (lfsr_C_1), .S0 (test_mode)) ;
    dff test_input_reg_BP2_1 (.Q (lfsr_C_1), .QB (\$dummy [20]), .D (
        test_input_lfsr_signal_1), .CLK (CLK)) ;
    aoi32 ix2596 (.Y (nx2595), .A0 (nx5448), .A1 (nx5464), .A2 (mac_unit_tempP_0
          ), .B0 (Cin), .B1 (nx1937)) ;
    nor02ii ix4315 (.Y (mac_output[2]), .A0 (RST), .A1 (nx4310)) ;
    nor02 ix4311 (.Y (nx4310), .A0 (RST), .A1 (nx2601)) ;
    xnor2 ix2602 (.Y (nx2601), .A0 (nx2603), .A1 (nx2609)) ;
    xnor2 ix2604 (.Y (nx2603), .A0 (mac_unit_tempP_2), .A1 (nx3692)) ;
    dffr mac_unit_MR_reg_Q_2 (.Q (mac_unit_tempP_2), .QB (\$dummy [21]), .D (
         nx3680), .CLK (CLK), .R (RST)) ;
    mux21 ix2610 (.Y (nx2609), .A0 (nx2565), .A1 (nx2595), .S0 (nx1935)) ;
    aoi21 ix3693 (.Y (nx3692), .A0 (nx2613), .A1 (nx2621), .B0 (nx688)) ;
    mux21 ix529 (.Y (nx528), .A0 (B[2]), .A1 (lfsr_C_13), .S0 (test_mode)) ;
    dff test_input_reg_BP2_13 (.Q (lfsr_C_13), .QB (\$dummy [22]), .D (
        test_input_lfsr_signal_13), .CLK (CLK)) ;
    xnor2 ix2622 (.Y (nx2621), .A0 (nx2567), .A1 (nx2623)) ;
    xnor2 ix2624 (.Y (nx2623), .A0 (nx2625), .A1 (nx2627)) ;
    nand02 ix2628 (.Y (nx2627), .A0 (nx5448), .A1 (nx410)) ;
    mux21 ix411 (.Y (nx410), .A0 (C[2]), .A1 (lfsr_C_2), .S0 (test_mode)) ;
    dff test_input_reg_BP2_2 (.Q (lfsr_C_2), .QB (\$dummy [23]), .D (
        test_input_lfsr_signal_2), .CLK (CLK)) ;
    nor03 ix689 (.Y (nx688), .A0 (nx2621), .A1 (nx5536), .A2 (nx2635)) ;
    nor02ii ix4323 (.Y (mac_output[3]), .A0 (RST), .A1 (nx4318)) ;
    nor02 ix4319 (.Y (nx4318), .A0 (RST), .A1 (nx2643)) ;
    xnor2 ix2644 (.Y (nx2643), .A0 (nx2645), .A1 (nx2651)) ;
    xnor2 ix2646 (.Y (nx2645), .A0 (mac_unit_tempP_3), .A1 (nx3716)) ;
    dffr mac_unit_MR_reg_Q_3 (.Q (mac_unit_tempP_3), .QB (\$dummy [24]), .D (
         nx3704), .CLK (CLK), .R (RST)) ;
    aoi22 ix2652 (.Y (nx2651), .A0 (nx3692), .A1 (mac_unit_tempP_2), .B0 (nx1933
          ), .B1 (nx3678)) ;
    aoi21 ix3717 (.Y (nx3716), .A0 (nx2661), .A1 (nx2668), .B0 (nx910)) ;
    mux21 ix757 (.Y (nx756), .A0 (B[3]), .A1 (lfsr_C_12), .S0 (test_mode)) ;
    dff test_input_reg_BP2_12 (.Q (lfsr_C_12), .QB (\$dummy [25]), .D (
        test_input_lfsr_signal_12), .CLK (CLK)) ;
    xnor2 ix2670 (.Y (nx2668), .A0 (nx688), .A1 (nx678)) ;
    xnor2 ix679 (.Y (nx678), .A0 (nx2673), .A1 (nx674)) ;
    xnor2 ix675 (.Y (nx674), .A0 (nx464), .A1 (nx2679)) ;
    aoi21 ix465 (.Y (nx464), .A0 (nx2439), .A1 (nx2627), .B0 (nx2625)) ;
    xnor2 ix2680 (.Y (nx2679), .A0 (nx2681), .A1 (nx2683)) ;
    nand02 ix2682 (.Y (nx2681), .A0 (nx5456), .A1 (nx410)) ;
    nand02 ix2684 (.Y (nx2683), .A0 (nx5448), .A1 (nx386)) ;
    mux21 ix387 (.Y (nx386), .A0 (C[3]), .A1 (lfsr_C_3), .S0 (test_mode)) ;
    dff test_input_reg_BP2_3 (.Q (lfsr_C_3), .QB (\$dummy [26]), .D (
        test_input_lfsr_signal_3), .CLK (CLK)) ;
    nor03 ix911 (.Y (nx910), .A0 (nx2668), .A1 (nx5536), .A2 (nx2691)) ;
    nor02ii ix4331 (.Y (mac_output[4]), .A0 (RST), .A1 (nx4326)) ;
    nor02 ix4327 (.Y (nx4326), .A0 (RST), .A1 (nx2699)) ;
    xnor2 ix2700 (.Y (nx2699), .A0 (nx2701), .A1 (nx2707)) ;
    xnor2 ix2702 (.Y (nx2701), .A0 (mac_unit_tempP_4), .A1 (nx3740)) ;
    dffr mac_unit_MR_reg_Q_4 (.Q (mac_unit_tempP_4), .QB (\$dummy [27]), .D (
         nx3728), .CLK (CLK), .R (RST)) ;
    aoi22 ix2708 (.Y (nx2707), .A0 (nx3716), .A1 (mac_unit_tempP_3), .B0 (nx1932
          ), .B1 (nx3702)) ;
    aoi21 ix3741 (.Y (nx3740), .A0 (nx2717), .A1 (nx2725), .B0 (nx1132)) ;
    mux21 ix979 (.Y (nx978), .A0 (B[4]), .A1 (lfsr_C_11), .S0 (test_mode)) ;
    dff test_input_reg_BP2_11 (.Q (lfsr_C_11), .QB (\$dummy [28]), .D (
        test_input_lfsr_signal_11), .CLK (CLK)) ;
    xnor2 ix2726 (.Y (nx2725), .A0 (nx910), .A1 (nx900)) ;
    xnor2 ix901 (.Y (nx900), .A0 (nx2729), .A1 (nx896)) ;
    xnor2 ix897 (.Y (nx896), .A0 (nx692), .A1 (nx2735)) ;
    mux21 ix693 (.Y (nx692), .A0 (nx674), .A1 (nx688), .S0 (nx678)) ;
    xnor2 ix2736 (.Y (nx2735), .A0 (nx2737), .A1 (nx2739)) ;
    nand02 ix2738 (.Y (nx2737), .A0 (nx5468), .A1 (nx410)) ;
    xnor2 ix2740 (.Y (nx2739), .A0 (nx2741), .A1 (nx2745)) ;
    mux21 ix2742 (.Y (nx2741), .A0 (nx2743), .A1 (nx2683), .S0 (nx2679)) ;
    xnor2 ix2746 (.Y (nx2745), .A0 (nx2747), .A1 (nx2749)) ;
    nand02 ix2748 (.Y (nx2747), .A0 (nx5456), .A1 (nx386)) ;
    nand02 ix2750 (.Y (nx2749), .A0 (nx5448), .A1 (nx362)) ;
    mux21 ix363 (.Y (nx362), .A0 (C[4]), .A1 (lfsr_C_4), .S0 (test_mode)) ;
    dff test_input_reg_BP2_4 (.Q (lfsr_C_4), .QB (\$dummy [29]), .D (
        test_input_lfsr_signal_4), .CLK (CLK)) ;
    nor03 ix1133 (.Y (nx1132), .A0 (nx2725), .A1 (nx5536), .A2 (nx2757)) ;
    nor02ii ix4339 (.Y (mac_output[5]), .A0 (RST), .A1 (nx4334)) ;
    nor02 ix4335 (.Y (nx4334), .A0 (RST), .A1 (nx2765)) ;
    xnor2 ix2766 (.Y (nx2765), .A0 (nx2767), .A1 (nx2773)) ;
    xnor2 ix2768 (.Y (nx2767), .A0 (mac_unit_tempP_5), .A1 (nx3764)) ;
    dffr mac_unit_MR_reg_Q_5 (.Q (mac_unit_tempP_5), .QB (\$dummy [30]), .D (
         nx3752), .CLK (CLK), .R (RST)) ;
    aoi22 ix2774 (.Y (nx2773), .A0 (nx3740), .A1 (mac_unit_tempP_4), .B0 (nx1931
          ), .B1 (nx3726)) ;
    aoi21 ix3765 (.Y (nx3764), .A0 (nx2783), .A1 (nx2790), .B0 (nx1354)) ;
    mux21 ix1201 (.Y (nx1200), .A0 (B[5]), .A1 (lfsr_C_10), .S0 (test_mode)) ;
    dff test_input_reg_BP2_10 (.Q (lfsr_C_10), .QB (\$dummy [31]), .D (
        test_input_lfsr_signal_10), .CLK (CLK)) ;
    xnor2 ix2792 (.Y (nx2790), .A0 (nx1132), .A1 (nx1122)) ;
    xnor2 ix1123 (.Y (nx1122), .A0 (nx2795), .A1 (nx1118)) ;
    xnor2 ix1119 (.Y (nx1118), .A0 (nx914), .A1 (nx2801)) ;
    mux21 ix915 (.Y (nx914), .A0 (nx896), .A1 (nx910), .S0 (nx900)) ;
    xnor2 ix2802 (.Y (nx2801), .A0 (nx2803), .A1 (nx2805)) ;
    nand02 ix2804 (.Y (nx2803), .A0 (nx410), .A1 (nx5472)) ;
    xnor2 ix2806 (.Y (nx2805), .A0 (nx2807), .A1 (nx2811)) ;
    mux21 ix2808 (.Y (nx2807), .A0 (nx2809), .A1 (nx2739), .S0 (nx2735)) ;
    xnor2 ix2812 (.Y (nx2811), .A0 (nx2813), .A1 (nx2815)) ;
    nand02 ix2814 (.Y (nx2813), .A0 (nx5468), .A1 (nx386)) ;
    xnor2 ix2816 (.Y (nx2815), .A0 (nx2817), .A1 (nx2819)) ;
    mux21 ix2818 (.Y (nx2817), .A0 (nx2741), .A1 (nx2749), .S0 (nx2745)) ;
    xnor2 ix2820 (.Y (nx2819), .A0 (nx2821), .A1 (nx2823)) ;
    nand02 ix2822 (.Y (nx2821), .A0 (nx5456), .A1 (nx362)) ;
    nand02 ix2824 (.Y (nx2823), .A0 (nx5448), .A1 (nx338)) ;
    mux21 ix339 (.Y (nx338), .A0 (C[5]), .A1 (lfsr_C_5), .S0 (test_mode)) ;
    dff test_input_reg_BP2_5 (.Q (lfsr_C_5), .QB (\$dummy [32]), .D (
        test_input_lfsr_signal_5), .CLK (CLK)) ;
    nor03 ix1355 (.Y (nx1354), .A0 (nx2790), .A1 (nx5536), .A2 (nx2831)) ;
    nor02ii ix4347 (.Y (mac_output[6]), .A0 (RST), .A1 (nx4342)) ;
    nor02 ix4343 (.Y (nx4342), .A0 (RST), .A1 (nx2839)) ;
    xnor2 ix2840 (.Y (nx2839), .A0 (nx2841), .A1 (nx2847)) ;
    xnor2 ix2842 (.Y (nx2841), .A0 (mac_unit_tempP_6), .A1 (nx3788)) ;
    dffr mac_unit_MR_reg_Q_6 (.Q (mac_unit_tempP_6), .QB (\$dummy [33]), .D (
         nx3776), .CLK (CLK), .R (RST)) ;
    aoi22 ix2848 (.Y (nx2847), .A0 (nx3764), .A1 (mac_unit_tempP_5), .B0 (nx1929
          ), .B1 (nx3750)) ;
    aoi21 ix3789 (.Y (nx3788), .A0 (nx2857), .A1 (nx2865), .B0 (nx1576)) ;
    mux21 ix1423 (.Y (nx1422), .A0 (B[6]), .A1 (lfsr_C_9), .S0 (test_mode)) ;
    dff test_input_reg_BP2_9 (.Q (lfsr_C_9), .QB (\$dummy [34]), .D (
        test_input_lfsr_signal_9), .CLK (CLK)) ;
    xnor2 ix2866 (.Y (nx2865), .A0 (nx1354), .A1 (nx1344)) ;
    xnor2 ix1345 (.Y (nx1344), .A0 (nx2869), .A1 (nx1340)) ;
    xnor2 ix1341 (.Y (nx1340), .A0 (nx1136), .A1 (nx2875)) ;
    mux21 ix1137 (.Y (nx1136), .A0 (nx1118), .A1 (nx1132), .S0 (nx1122)) ;
    xnor2 ix2876 (.Y (nx2875), .A0 (nx2877), .A1 (nx2879)) ;
    nand02 ix2878 (.Y (nx2877), .A0 (nx410), .A1 (nx5476)) ;
    xnor2 ix2880 (.Y (nx2879), .A0 (nx2881), .A1 (nx2885)) ;
    mux21 ix2882 (.Y (nx2881), .A0 (nx2883), .A1 (nx2805), .S0 (nx2801)) ;
    xnor2 ix2886 (.Y (nx2885), .A0 (nx2887), .A1 (nx2889)) ;
    nand02 ix2888 (.Y (nx2887), .A0 (nx5472), .A1 (nx386)) ;
    xnor2 ix2890 (.Y (nx2889), .A0 (nx2891), .A1 (nx2893)) ;
    mux21 ix2892 (.Y (nx2891), .A0 (nx2807), .A1 (nx2815), .S0 (nx2811)) ;
    xnor2 ix2894 (.Y (nx2893), .A0 (nx2895), .A1 (nx2897)) ;
    nand02 ix2896 (.Y (nx2895), .A0 (nx5468), .A1 (nx362)) ;
    xnor2 ix2898 (.Y (nx2897), .A0 (nx2899), .A1 (nx2901)) ;
    mux21 ix2900 (.Y (nx2899), .A0 (nx2817), .A1 (nx2823), .S0 (nx2819)) ;
    xnor2 ix2902 (.Y (nx2901), .A0 (nx2903), .A1 (nx2905)) ;
    nand02 ix2904 (.Y (nx2903), .A0 (nx5456), .A1 (nx338)) ;
    nand02 ix2906 (.Y (nx2905), .A0 (nx5448), .A1 (nx314)) ;
    mux21 ix315 (.Y (nx314), .A0 (C[6]), .A1 (lfsr_C_6), .S0 (test_mode)) ;
    dff test_input_reg_BP2_6 (.Q (lfsr_C_6), .QB (\$dummy [35]), .D (
        test_input_lfsr_signal_6), .CLK (CLK)) ;
    nor03 ix1577 (.Y (nx1576), .A0 (nx2865), .A1 (nx5536), .A2 (nx2913)) ;
    nor02ii ix4355 (.Y (mac_output[7]), .A0 (RST), .A1 (nx4350)) ;
    nor02 ix4351 (.Y (nx4350), .A0 (RST), .A1 (nx2921)) ;
    xnor2 ix2922 (.Y (nx2921), .A0 (nx2923), .A1 (nx2929)) ;
    xnor2 ix2924 (.Y (nx2923), .A0 (mac_unit_tempP_7), .A1 (nx3812)) ;
    dffr mac_unit_MR_reg_Q_7 (.Q (mac_unit_tempP_7), .QB (\$dummy [36]), .D (
         nx3800), .CLK (CLK), .R (RST)) ;
    aoi22 ix2930 (.Y (nx2929), .A0 (nx3788), .A1 (mac_unit_tempP_6), .B0 (nx1927
          ), .B1 (nx3774)) ;
    aoi21 ix3813 (.Y (nx3812), .A0 (nx2939), .A1 (nx2947), .B0 (nx1798)) ;
    mux21 ix1645 (.Y (nx1644), .A0 (B[7]), .A1 (lfsr_C_8), .S0 (test_mode)) ;
    dff test_input_reg_BP2_8 (.Q (lfsr_C_8), .QB (\$dummy [37]), .D (
        test_input_lfsr_signal_8), .CLK (CLK)) ;
    xnor2 ix2948 (.Y (nx2947), .A0 (nx1576), .A1 (nx1566)) ;
    xnor2 ix1567 (.Y (nx1566), .A0 (nx2951), .A1 (nx1562)) ;
    xnor2 ix1563 (.Y (nx1562), .A0 (nx1358), .A1 (nx2957)) ;
    mux21 ix1359 (.Y (nx1358), .A0 (nx1340), .A1 (nx1354), .S0 (nx1344)) ;
    xnor2 ix2958 (.Y (nx2957), .A0 (nx2959), .A1 (nx2961)) ;
    nand02 ix2960 (.Y (nx2959), .A0 (nx410), .A1 (nx5480)) ;
    xnor2 ix2962 (.Y (nx2961), .A0 (nx2963), .A1 (nx2967)) ;
    mux21 ix2964 (.Y (nx2963), .A0 (nx2965), .A1 (nx2879), .S0 (nx2875)) ;
    xnor2 ix2968 (.Y (nx2967), .A0 (nx2969), .A1 (nx2971)) ;
    nand02 ix2970 (.Y (nx2969), .A0 (nx386), .A1 (nx5476)) ;
    xnor2 ix2972 (.Y (nx2971), .A0 (nx2973), .A1 (nx2975)) ;
    mux21 ix2974 (.Y (nx2973), .A0 (nx2881), .A1 (nx2889), .S0 (nx2885)) ;
    xnor2 ix2976 (.Y (nx2975), .A0 (nx2977), .A1 (nx2979)) ;
    nand02 ix2978 (.Y (nx2977), .A0 (nx5472), .A1 (nx362)) ;
    xnor2 ix2980 (.Y (nx2979), .A0 (nx2981), .A1 (nx2983)) ;
    mux21 ix2982 (.Y (nx2981), .A0 (nx2891), .A1 (nx2897), .S0 (nx2893)) ;
    xnor2 ix2984 (.Y (nx2983), .A0 (nx2985), .A1 (nx2987)) ;
    nand02 ix2986 (.Y (nx2985), .A0 (nx5468), .A1 (nx338)) ;
    xnor2 ix2988 (.Y (nx2987), .A0 (nx2989), .A1 (nx2991)) ;
    mux21 ix2990 (.Y (nx2989), .A0 (nx2899), .A1 (nx2905), .S0 (nx2901)) ;
    xnor2 ix2992 (.Y (nx2991), .A0 (nx2993), .A1 (nx2995)) ;
    nand02 ix2994 (.Y (nx2993), .A0 (nx5456), .A1 (nx314)) ;
    nand02 ix2996 (.Y (nx2995), .A0 (nx5448), .A1 (nx290)) ;
    mux21 ix291 (.Y (nx290), .A0 (C[7]), .A1 (lfsr_C_7), .S0 (test_mode)) ;
    dff test_input_reg_BP2_7 (.Q (lfsr_C_7), .QB (\$dummy [38]), .D (
        test_input_lfsr_signal_7), .CLK (CLK)) ;
    nor03 ix1799 (.Y (nx1798), .A0 (nx2947), .A1 (nx5536), .A2 (nx3003)) ;
    nor02ii ix4363 (.Y (mac_output[8]), .A0 (RST), .A1 (nx4358)) ;
    nor02 ix4359 (.Y (nx4358), .A0 (RST), .A1 (nx3011)) ;
    xnor2 ix3012 (.Y (nx3011), .A0 (nx3013), .A1 (nx3019)) ;
    xnor2 ix3014 (.Y (nx3013), .A0 (mac_unit_tempP_8), .A1 (nx3836)) ;
    dffr mac_unit_MR_reg_Q_8 (.Q (mac_unit_tempP_8), .QB (\$dummy [39]), .D (
         nx3824), .CLK (CLK), .R (RST)) ;
    aoi22 ix3020 (.Y (nx3019), .A0 (nx3812), .A1 (mac_unit_tempP_7), .B0 (nx1925
          ), .B1 (nx3798)) ;
    aoi21 ix3837 (.Y (nx3836), .A0 (nx3029), .A1 (nx3033), .B0 (nx2020)) ;
    mux21 ix1867 (.Y (nx1866), .A0 (B[8]), .A1 (lfsr_C_7), .S0 (test_mode)) ;
    xnor2 ix3034 (.Y (nx3033), .A0 (nx1798), .A1 (nx1788)) ;
    xnor2 ix1789 (.Y (nx1788), .A0 (nx3037), .A1 (nx1784)) ;
    xnor2 ix1785 (.Y (nx1784), .A0 (nx1580), .A1 (nx3043)) ;
    mux21 ix1581 (.Y (nx1580), .A0 (nx1562), .A1 (nx1576), .S0 (nx1566)) ;
    xnor2 ix3044 (.Y (nx3043), .A0 (nx3045), .A1 (nx3047)) ;
    nand02 ix3046 (.Y (nx3045), .A0 (nx410), .A1 (nx5484)) ;
    xnor2 ix3048 (.Y (nx3047), .A0 (nx3049), .A1 (nx3053)) ;
    mux21 ix3050 (.Y (nx3049), .A0 (nx3051), .A1 (nx2961), .S0 (nx2957)) ;
    xnor2 ix3054 (.Y (nx3053), .A0 (nx3055), .A1 (nx3057)) ;
    nand02 ix3056 (.Y (nx3055), .A0 (nx386), .A1 (nx5480)) ;
    xnor2 ix3058 (.Y (nx3057), .A0 (nx3059), .A1 (nx3061)) ;
    mux21 ix3060 (.Y (nx3059), .A0 (nx2963), .A1 (nx2971), .S0 (nx2967)) ;
    xnor2 ix3062 (.Y (nx3061), .A0 (nx3063), .A1 (nx3065)) ;
    nand02 ix3064 (.Y (nx3063), .A0 (nx5476), .A1 (nx362)) ;
    xnor2 ix3066 (.Y (nx3065), .A0 (nx3067), .A1 (nx3069)) ;
    mux21 ix3068 (.Y (nx3067), .A0 (nx2973), .A1 (nx2979), .S0 (nx2975)) ;
    xnor2 ix3070 (.Y (nx3069), .A0 (nx3071), .A1 (nx3073)) ;
    nand02 ix3072 (.Y (nx3071), .A0 (nx5472), .A1 (nx338)) ;
    xnor2 ix3074 (.Y (nx3073), .A0 (nx3075), .A1 (nx3077)) ;
    mux21 ix3076 (.Y (nx3075), .A0 (nx2981), .A1 (nx2987), .S0 (nx2983)) ;
    xnor2 ix3078 (.Y (nx3077), .A0 (nx3079), .A1 (nx3081)) ;
    nand02 ix3080 (.Y (nx3079), .A0 (nx5468), .A1 (nx314)) ;
    xnor2 ix3082 (.Y (nx3081), .A0 (nx3083), .A1 (nx3085)) ;
    mux21 ix3084 (.Y (nx3083), .A0 (nx2989), .A1 (nx2995), .S0 (nx2991)) ;
    xnor2 ix3086 (.Y (nx3085), .A0 (nx3087), .A1 (nx3089)) ;
    nand02 ix3088 (.Y (nx3087), .A0 (nx5456), .A1 (nx290)) ;
    nand02 ix3090 (.Y (nx3089), .A0 (nx5448), .A1 (nx266)) ;
    mux21 ix267 (.Y (nx266), .A0 (C[8]), .A1 (lfsr_C_8), .S0 (test_mode)) ;
    nor03 ix2021 (.Y (nx2020), .A0 (nx3033), .A1 (nx5536), .A2 (nx3095)) ;
    nor02ii ix4371 (.Y (mac_output[9]), .A0 (RST), .A1 (nx4366)) ;
    nor02 ix4367 (.Y (nx4366), .A0 (RST), .A1 (nx3103)) ;
    xnor2 ix3104 (.Y (nx3103), .A0 (nx3105), .A1 (nx3111)) ;
    xnor2 ix3106 (.Y (nx3105), .A0 (mac_unit_tempP_9), .A1 (nx3860)) ;
    dffr mac_unit_MR_reg_Q_9 (.Q (mac_unit_tempP_9), .QB (\$dummy [40]), .D (
         nx3848), .CLK (CLK), .R (RST)) ;
    aoi22 ix3112 (.Y (nx3111), .A0 (nx3836), .A1 (mac_unit_tempP_8), .B0 (nx1923
          ), .B1 (nx3822)) ;
    aoi21 ix3861 (.Y (nx3860), .A0 (nx3121), .A1 (nx3125), .B0 (nx2242)) ;
    mux21 ix2089 (.Y (nx2088), .A0 (B[9]), .A1 (lfsr_C_6), .S0 (test_mode)) ;
    xnor2 ix3126 (.Y (nx3125), .A0 (nx2020), .A1 (nx2010)) ;
    xnor2 ix2011 (.Y (nx2010), .A0 (nx3129), .A1 (nx2006)) ;
    xnor2 ix2007 (.Y (nx2006), .A0 (nx1802), .A1 (nx3135)) ;
    mux21 ix1803 (.Y (nx1802), .A0 (nx1784), .A1 (nx1798), .S0 (nx1788)) ;
    xnor2 ix3136 (.Y (nx3135), .A0 (nx3137), .A1 (nx3139)) ;
    nand02 ix3138 (.Y (nx3137), .A0 (nx410), .A1 (nx5488)) ;
    xnor2 ix3140 (.Y (nx3139), .A0 (nx3141), .A1 (nx3145)) ;
    mux21 ix3142 (.Y (nx3141), .A0 (nx3143), .A1 (nx3047), .S0 (nx3043)) ;
    xnor2 ix3146 (.Y (nx3145), .A0 (nx3147), .A1 (nx3149)) ;
    nand02 ix3148 (.Y (nx3147), .A0 (nx386), .A1 (nx5484)) ;
    xnor2 ix3150 (.Y (nx3149), .A0 (nx3151), .A1 (nx3153)) ;
    mux21 ix3152 (.Y (nx3151), .A0 (nx3049), .A1 (nx3057), .S0 (nx3053)) ;
    xnor2 ix3154 (.Y (nx3153), .A0 (nx3155), .A1 (nx3157)) ;
    nand02 ix3156 (.Y (nx3155), .A0 (nx362), .A1 (nx5480)) ;
    xnor2 ix3158 (.Y (nx3157), .A0 (nx3159), .A1 (nx3161)) ;
    mux21 ix3160 (.Y (nx3159), .A0 (nx3059), .A1 (nx3065), .S0 (nx3061)) ;
    xnor2 ix3162 (.Y (nx3161), .A0 (nx3163), .A1 (nx3165)) ;
    nand02 ix3164 (.Y (nx3163), .A0 (nx5476), .A1 (nx338)) ;
    xnor2 ix3166 (.Y (nx3165), .A0 (nx3167), .A1 (nx3169)) ;
    mux21 ix3168 (.Y (nx3167), .A0 (nx3067), .A1 (nx3073), .S0 (nx3069)) ;
    xnor2 ix3170 (.Y (nx3169), .A0 (nx3171), .A1 (nx3173)) ;
    nand02 ix3172 (.Y (nx3171), .A0 (nx5472), .A1 (nx314)) ;
    xnor2 ix3174 (.Y (nx3173), .A0 (nx3175), .A1 (nx3177)) ;
    mux21 ix3176 (.Y (nx3175), .A0 (nx3075), .A1 (nx3081), .S0 (nx3077)) ;
    xnor2 ix3178 (.Y (nx3177), .A0 (nx3179), .A1 (nx3181)) ;
    nand02 ix3180 (.Y (nx3179), .A0 (nx5468), .A1 (nx290)) ;
    xnor2 ix3182 (.Y (nx3181), .A0 (nx3183), .A1 (nx3185)) ;
    mux21 ix3184 (.Y (nx3183), .A0 (nx3083), .A1 (nx3089), .S0 (nx3085)) ;
    xnor2 ix3186 (.Y (nx3185), .A0 (nx3187), .A1 (nx3189)) ;
    nand02 ix3188 (.Y (nx3187), .A0 (nx5456), .A1 (nx266)) ;
    nand02 ix3190 (.Y (nx3189), .A0 (nx5448), .A1 (nx242)) ;
    mux21 ix243 (.Y (nx242), .A0 (C[9]), .A1 (lfsr_C_9), .S0 (test_mode)) ;
    nor03 ix2243 (.Y (nx2242), .A0 (nx3125), .A1 (nx5536), .A2 (nx3195)) ;
    nor02ii ix4379 (.Y (mac_output[10]), .A0 (RST), .A1 (nx4374)) ;
    nor02 ix4375 (.Y (nx4374), .A0 (RST), .A1 (nx3203)) ;
    xnor2 ix3204 (.Y (nx3203), .A0 (nx3205), .A1 (nx3211)) ;
    xnor2 ix3206 (.Y (nx3205), .A0 (mac_unit_tempP_10), .A1 (nx3884)) ;
    dffr mac_unit_MR_reg_Q_10 (.Q (mac_unit_tempP_10), .QB (\$dummy [41]), .D (
         nx3872), .CLK (CLK), .R (RST)) ;
    aoi22 ix3212 (.Y (nx3211), .A0 (nx3860), .A1 (mac_unit_tempP_9), .B0 (nx1922
          ), .B1 (nx3846)) ;
    aoi21 ix3885 (.Y (nx3884), .A0 (nx3221), .A1 (nx3225), .B0 (nx2464)) ;
    mux21 ix2311 (.Y (nx2310), .A0 (B[10]), .A1 (lfsr_C_5), .S0 (test_mode)) ;
    xnor2 ix3226 (.Y (nx3225), .A0 (nx2242), .A1 (nx2232)) ;
    xnor2 ix2233 (.Y (nx2232), .A0 (nx3229), .A1 (nx2228)) ;
    xnor2 ix2229 (.Y (nx2228), .A0 (nx2024), .A1 (nx3235)) ;
    mux21 ix2025 (.Y (nx2024), .A0 (nx2006), .A1 (nx2020), .S0 (nx2010)) ;
    xnor2 ix3236 (.Y (nx3235), .A0 (nx3237), .A1 (nx3239)) ;
    nand02 ix3238 (.Y (nx3237), .A0 (nx410), .A1 (nx5492)) ;
    xnor2 ix3240 (.Y (nx3239), .A0 (nx3241), .A1 (nx3245)) ;
    mux21 ix3242 (.Y (nx3241), .A0 (nx3243), .A1 (nx3139), .S0 (nx3135)) ;
    xnor2 ix3246 (.Y (nx3245), .A0 (nx3247), .A1 (nx3249)) ;
    nand02 ix3248 (.Y (nx3247), .A0 (nx386), .A1 (nx5488)) ;
    xnor2 ix3250 (.Y (nx3249), .A0 (nx3251), .A1 (nx3253)) ;
    mux21 ix3252 (.Y (nx3251), .A0 (nx3141), .A1 (nx3149), .S0 (nx3145)) ;
    xnor2 ix3254 (.Y (nx3253), .A0 (nx3255), .A1 (nx3257)) ;
    nand02 ix3256 (.Y (nx3255), .A0 (nx362), .A1 (nx5484)) ;
    xnor2 ix3258 (.Y (nx3257), .A0 (nx3259), .A1 (nx3261)) ;
    mux21 ix3260 (.Y (nx3259), .A0 (nx3151), .A1 (nx3157), .S0 (nx3153)) ;
    xnor2 ix3262 (.Y (nx3261), .A0 (nx3263), .A1 (nx3265)) ;
    nand02 ix3264 (.Y (nx3263), .A0 (nx5480), .A1 (nx338)) ;
    xnor2 ix3266 (.Y (nx3265), .A0 (nx3267), .A1 (nx3269)) ;
    mux21 ix3268 (.Y (nx3267), .A0 (nx3159), .A1 (nx3165), .S0 (nx3161)) ;
    xnor2 ix3270 (.Y (nx3269), .A0 (nx3271), .A1 (nx3273)) ;
    nand02 ix3272 (.Y (nx3271), .A0 (nx5476), .A1 (nx314)) ;
    xnor2 ix3274 (.Y (nx3273), .A0 (nx3275), .A1 (nx3277)) ;
    mux21 ix3276 (.Y (nx3275), .A0 (nx3167), .A1 (nx3173), .S0 (nx3169)) ;
    xnor2 ix3278 (.Y (nx3277), .A0 (nx3279), .A1 (nx3281)) ;
    nand02 ix3280 (.Y (nx3279), .A0 (nx5472), .A1 (nx290)) ;
    xnor2 ix3282 (.Y (nx3281), .A0 (nx3283), .A1 (nx3285)) ;
    mux21 ix3284 (.Y (nx3283), .A0 (nx3175), .A1 (nx3181), .S0 (nx3177)) ;
    xnor2 ix3286 (.Y (nx3285), .A0 (nx3287), .A1 (nx3289)) ;
    nand02 ix3288 (.Y (nx3287), .A0 (nx5468), .A1 (nx266)) ;
    xnor2 ix3290 (.Y (nx3289), .A0 (nx3291), .A1 (nx3293)) ;
    mux21 ix3292 (.Y (nx3291), .A0 (nx3183), .A1 (nx3189), .S0 (nx3185)) ;
    xnor2 ix3294 (.Y (nx3293), .A0 (nx3295), .A1 (nx3297)) ;
    nand02 ix3296 (.Y (nx3295), .A0 (nx5456), .A1 (nx242)) ;
    nand02 ix3298 (.Y (nx3297), .A0 (nx5448), .A1 (nx218)) ;
    mux21 ix219 (.Y (nx218), .A0 (C[10]), .A1 (lfsr_C_10), .S0 (test_mode)) ;
    nor03 ix2465 (.Y (nx2464), .A0 (nx3225), .A1 (nx5536), .A2 (nx3303)) ;
    nor02ii ix4387 (.Y (mac_output[11]), .A0 (RST), .A1 (nx4382)) ;
    nor02 ix4383 (.Y (nx4382), .A0 (RST), .A1 (nx3311)) ;
    xnor2 ix3312 (.Y (nx3311), .A0 (nx3313), .A1 (nx3319)) ;
    xnor2 ix3314 (.Y (nx3313), .A0 (mac_unit_tempP_11), .A1 (nx3908)) ;
    dffr mac_unit_MR_reg_Q_11 (.Q (mac_unit_tempP_11), .QB (\$dummy [42]), .D (
         nx3896), .CLK (CLK), .R (RST)) ;
    aoi22 ix3320 (.Y (nx3319), .A0 (nx3884), .A1 (mac_unit_tempP_10), .B0 (
          nx1921), .B1 (nx3870)) ;
    aoi21 ix3909 (.Y (nx3908), .A0 (nx3329), .A1 (nx3333), .B0 (nx2686)) ;
    mux21 ix2533 (.Y (nx2532), .A0 (B[11]), .A1 (lfsr_C_4), .S0 (test_mode)) ;
    xnor2 ix3334 (.Y (nx3333), .A0 (nx2464), .A1 (nx2454)) ;
    xnor2 ix2455 (.Y (nx2454), .A0 (nx3337), .A1 (nx2450)) ;
    xnor2 ix2451 (.Y (nx2450), .A0 (nx2246), .A1 (nx3343)) ;
    mux21 ix2247 (.Y (nx2246), .A0 (nx2228), .A1 (nx2242), .S0 (nx2232)) ;
    xnor2 ix3344 (.Y (nx3343), .A0 (nx3345), .A1 (nx3347)) ;
    nand02 ix3346 (.Y (nx3345), .A0 (nx410), .A1 (nx5496)) ;
    xnor2 ix3348 (.Y (nx3347), .A0 (nx3349), .A1 (nx3353)) ;
    mux21 ix3350 (.Y (nx3349), .A0 (nx3351), .A1 (nx3239), .S0 (nx3235)) ;
    xnor2 ix3354 (.Y (nx3353), .A0 (nx3355), .A1 (nx3357)) ;
    nand02 ix3356 (.Y (nx3355), .A0 (nx386), .A1 (nx5492)) ;
    xnor2 ix3358 (.Y (nx3357), .A0 (nx3359), .A1 (nx3361)) ;
    mux21 ix3360 (.Y (nx3359), .A0 (nx3241), .A1 (nx3249), .S0 (nx3245)) ;
    xnor2 ix3362 (.Y (nx3361), .A0 (nx3363), .A1 (nx3365)) ;
    nand02 ix3364 (.Y (nx3363), .A0 (nx362), .A1 (nx5488)) ;
    xnor2 ix3366 (.Y (nx3365), .A0 (nx3367), .A1 (nx3369)) ;
    mux21 ix3368 (.Y (nx3367), .A0 (nx3251), .A1 (nx3257), .S0 (nx3253)) ;
    xnor2 ix3370 (.Y (nx3369), .A0 (nx3371), .A1 (nx3373)) ;
    nand02 ix3372 (.Y (nx3371), .A0 (nx338), .A1 (nx5484)) ;
    xnor2 ix3374 (.Y (nx3373), .A0 (nx3375), .A1 (nx3377)) ;
    mux21 ix3376 (.Y (nx3375), .A0 (nx3259), .A1 (nx3265), .S0 (nx3261)) ;
    xnor2 ix3378 (.Y (nx3377), .A0 (nx3379), .A1 (nx3381)) ;
    nand02 ix3380 (.Y (nx3379), .A0 (nx5480), .A1 (nx314)) ;
    xnor2 ix3382 (.Y (nx3381), .A0 (nx3383), .A1 (nx3385)) ;
    mux21 ix3384 (.Y (nx3383), .A0 (nx3267), .A1 (nx3273), .S0 (nx3269)) ;
    xnor2 ix3386 (.Y (nx3385), .A0 (nx3387), .A1 (nx3389)) ;
    nand02 ix3388 (.Y (nx3387), .A0 (nx5476), .A1 (nx290)) ;
    xnor2 ix3390 (.Y (nx3389), .A0 (nx3391), .A1 (nx3393)) ;
    mux21 ix3392 (.Y (nx3391), .A0 (nx3275), .A1 (nx3281), .S0 (nx3277)) ;
    xnor2 ix3394 (.Y (nx3393), .A0 (nx3395), .A1 (nx3397)) ;
    nand02 ix3396 (.Y (nx3395), .A0 (nx5472), .A1 (nx266)) ;
    xnor2 ix3398 (.Y (nx3397), .A0 (nx3399), .A1 (nx3401)) ;
    mux21 ix3400 (.Y (nx3399), .A0 (nx3283), .A1 (nx3289), .S0 (nx3285)) ;
    xnor2 ix3402 (.Y (nx3401), .A0 (nx3403), .A1 (nx3405)) ;
    nand02 ix3404 (.Y (nx3403), .A0 (nx5468), .A1 (nx242)) ;
    xnor2 ix3406 (.Y (nx3405), .A0 (nx3407), .A1 (nx3409)) ;
    mux21 ix3408 (.Y (nx3407), .A0 (nx3291), .A1 (nx3297), .S0 (nx3293)) ;
    xnor2 ix3410 (.Y (nx3409), .A0 (nx3411), .A1 (nx3413)) ;
    nand02 ix3412 (.Y (nx3411), .A0 (nx5456), .A1 (nx218)) ;
    nand02 ix3414 (.Y (nx3413), .A0 (nx5448), .A1 (nx194)) ;
    mux21 ix195 (.Y (nx194), .A0 (C[11]), .A1 (lfsr_C_11), .S0 (test_mode)) ;
    nor03 ix2687 (.Y (nx2686), .A0 (nx3333), .A1 (nx5536), .A2 (nx3417)) ;
    nor02ii ix4395 (.Y (mac_output[12]), .A0 (RST), .A1 (nx4390)) ;
    nor02 ix4391 (.Y (nx4390), .A0 (RST), .A1 (nx3425)) ;
    xnor2 ix3426 (.Y (nx3425), .A0 (nx3427), .A1 (nx3433)) ;
    xnor2 ix3428 (.Y (nx3427), .A0 (mac_unit_tempP_12), .A1 (nx3932)) ;
    dffr mac_unit_MR_reg_Q_12 (.Q (mac_unit_tempP_12), .QB (\$dummy [43]), .D (
         nx3920), .CLK (CLK), .R (RST)) ;
    aoi22 ix3434 (.Y (nx3433), .A0 (nx3908), .A1 (mac_unit_tempP_11), .B0 (
          nx1919), .B1 (nx3894)) ;
    aoi21 ix3933 (.Y (nx3932), .A0 (nx3443), .A1 (nx3447), .B0 (nx2908)) ;
    mux21 ix2755 (.Y (nx2754), .A0 (B[12]), .A1 (lfsr_C_3), .S0 (test_mode)) ;
    xnor2 ix3448 (.Y (nx3447), .A0 (nx2686), .A1 (nx2676)) ;
    xnor2 ix2677 (.Y (nx2676), .A0 (nx3451), .A1 (nx2672)) ;
    xnor2 ix2673 (.Y (nx2672), .A0 (nx2468), .A1 (nx3457)) ;
    mux21 ix2469 (.Y (nx2468), .A0 (nx2450), .A1 (nx2464), .S0 (nx2454)) ;
    xnor2 ix3458 (.Y (nx3457), .A0 (nx3459), .A1 (nx3461)) ;
    nand02 ix3460 (.Y (nx3459), .A0 (nx410), .A1 (nx5500)) ;
    xnor2 ix3462 (.Y (nx3461), .A0 (nx3463), .A1 (nx3467)) ;
    mux21 ix3464 (.Y (nx3463), .A0 (nx3465), .A1 (nx3347), .S0 (nx3343)) ;
    xnor2 ix3468 (.Y (nx3467), .A0 (nx3469), .A1 (nx3471)) ;
    nand02 ix3470 (.Y (nx3469), .A0 (nx386), .A1 (nx5496)) ;
    xnor2 ix3472 (.Y (nx3471), .A0 (nx3473), .A1 (nx3475)) ;
    mux21 ix3474 (.Y (nx3473), .A0 (nx3349), .A1 (nx3357), .S0 (nx3353)) ;
    xnor2 ix3476 (.Y (nx3475), .A0 (nx3477), .A1 (nx3479)) ;
    nand02 ix3478 (.Y (nx3477), .A0 (nx362), .A1 (nx5492)) ;
    xnor2 ix3480 (.Y (nx3479), .A0 (nx3481), .A1 (nx3483)) ;
    mux21 ix3482 (.Y (nx3481), .A0 (nx3359), .A1 (nx3365), .S0 (nx3361)) ;
    xnor2 ix3484 (.Y (nx3483), .A0 (nx3485), .A1 (nx3487)) ;
    nand02 ix3486 (.Y (nx3485), .A0 (nx338), .A1 (nx5488)) ;
    xnor2 ix3488 (.Y (nx3487), .A0 (nx3489), .A1 (nx3491)) ;
    mux21 ix3490 (.Y (nx3489), .A0 (nx3367), .A1 (nx3373), .S0 (nx3369)) ;
    xnor2 ix3492 (.Y (nx3491), .A0 (nx3493), .A1 (nx3495)) ;
    nand02 ix3494 (.Y (nx3493), .A0 (nx5484), .A1 (nx314)) ;
    xnor2 ix3496 (.Y (nx3495), .A0 (nx3497), .A1 (nx3499)) ;
    mux21 ix3498 (.Y (nx3497), .A0 (nx3375), .A1 (nx3381), .S0 (nx3377)) ;
    xnor2 ix3500 (.Y (nx3499), .A0 (nx3501), .A1 (nx3503)) ;
    nand02 ix3502 (.Y (nx3501), .A0 (nx5480), .A1 (nx290)) ;
    xnor2 ix3504 (.Y (nx3503), .A0 (nx3505), .A1 (nx3507)) ;
    mux21 ix3506 (.Y (nx3505), .A0 (nx3383), .A1 (nx3389), .S0 (nx3385)) ;
    xnor2 ix3508 (.Y (nx3507), .A0 (nx3509), .A1 (nx3511)) ;
    nand02 ix3510 (.Y (nx3509), .A0 (nx5476), .A1 (nx266)) ;
    xnor2 ix3512 (.Y (nx3511), .A0 (nx3513), .A1 (nx3515)) ;
    mux21 ix3514 (.Y (nx3513), .A0 (nx3391), .A1 (nx3397), .S0 (nx3393)) ;
    xnor2 ix3516 (.Y (nx3515), .A0 (nx3517), .A1 (nx3519)) ;
    nand02 ix3518 (.Y (nx3517), .A0 (nx5472), .A1 (nx242)) ;
    xnor2 ix3520 (.Y (nx3519), .A0 (nx3521), .A1 (nx3523)) ;
    mux21 ix3522 (.Y (nx3521), .A0 (nx3399), .A1 (nx3405), .S0 (nx3401)) ;
    xnor2 ix3524 (.Y (nx3523), .A0 (nx3525), .A1 (nx3527)) ;
    nand02 ix3526 (.Y (nx3525), .A0 (nx5468), .A1 (nx218)) ;
    xnor2 ix3528 (.Y (nx3527), .A0 (nx3529), .A1 (nx3531)) ;
    mux21 ix3530 (.Y (nx3529), .A0 (nx3407), .A1 (nx3413), .S0 (nx3409)) ;
    xnor2 ix3532 (.Y (nx3531), .A0 (nx3533), .A1 (nx3535)) ;
    nand02 ix3534 (.Y (nx3533), .A0 (nx5456), .A1 (nx194)) ;
    nand02 ix3536 (.Y (nx3535), .A0 (nx5448), .A1 (nx170)) ;
    mux21 ix171 (.Y (nx170), .A0 (C[12]), .A1 (lfsr_C_12), .S0 (test_mode)) ;
    nor03 ix2909 (.Y (nx2908), .A0 (nx3447), .A1 (nx5536), .A2 (nx3541)) ;
    nor02ii ix4403 (.Y (mac_output[13]), .A0 (RST), .A1 (nx4398)) ;
    nor02 ix4399 (.Y (nx4398), .A0 (RST), .A1 (nx3549)) ;
    xnor2 ix3550 (.Y (nx3549), .A0 (nx3551), .A1 (nx3557)) ;
    xnor2 ix3552 (.Y (nx3551), .A0 (mac_unit_tempP_13), .A1 (nx3956)) ;
    dffr mac_unit_MR_reg_Q_13 (.Q (mac_unit_tempP_13), .QB (\$dummy [44]), .D (
         nx3944), .CLK (CLK), .R (RST)) ;
    aoi22 ix3558 (.Y (nx3557), .A0 (nx3932), .A1 (mac_unit_tempP_12), .B0 (
          nx1917), .B1 (nx3918)) ;
    aoi21 ix3957 (.Y (nx3956), .A0 (nx3567), .A1 (nx3571), .B0 (nx3130)) ;
    mux21 ix2977 (.Y (nx2976), .A0 (B[13]), .A1 (lfsr_C_2), .S0 (test_mode)) ;
    xnor2 ix3572 (.Y (nx3571), .A0 (nx2908), .A1 (nx2898)) ;
    xnor2 ix2899 (.Y (nx2898), .A0 (nx3575), .A1 (nx2894)) ;
    xnor2 ix2895 (.Y (nx2894), .A0 (nx2690), .A1 (nx3581)) ;
    mux21 ix2691 (.Y (nx2690), .A0 (nx2672), .A1 (nx2686), .S0 (nx2676)) ;
    xnor2 ix3582 (.Y (nx3581), .A0 (nx3583), .A1 (nx3585)) ;
    nand02 ix3584 (.Y (nx3583), .A0 (nx410), .A1 (nx5504)) ;
    xnor2 ix3586 (.Y (nx3585), .A0 (nx3587), .A1 (nx3591)) ;
    mux21 ix3588 (.Y (nx3587), .A0 (nx3589), .A1 (nx3461), .S0 (nx3457)) ;
    xnor2 ix3592 (.Y (nx3591), .A0 (nx3593), .A1 (nx3595)) ;
    nand02 ix3594 (.Y (nx3593), .A0 (nx386), .A1 (nx5500)) ;
    xnor2 ix3596 (.Y (nx3595), .A0 (nx3597), .A1 (nx3599)) ;
    mux21 ix3598 (.Y (nx3597), .A0 (nx3463), .A1 (nx3471), .S0 (nx3467)) ;
    xnor2 ix3600 (.Y (nx3599), .A0 (nx3601), .A1 (nx3603)) ;
    nand02 ix3602 (.Y (nx3601), .A0 (nx362), .A1 (nx5496)) ;
    xnor2 ix3604 (.Y (nx3603), .A0 (nx3605), .A1 (nx3607)) ;
    mux21 ix3606 (.Y (nx3605), .A0 (nx3473), .A1 (nx3479), .S0 (nx3475)) ;
    xnor2 ix3608 (.Y (nx3607), .A0 (nx3609), .A1 (nx3611)) ;
    nand02 ix3610 (.Y (nx3609), .A0 (nx338), .A1 (nx5492)) ;
    xnor2 ix3612 (.Y (nx3611), .A0 (nx3613), .A1 (nx3615)) ;
    mux21 ix3614 (.Y (nx3613), .A0 (nx3481), .A1 (nx3487), .S0 (nx3483)) ;
    xnor2 ix3616 (.Y (nx3615), .A0 (nx3617), .A1 (nx3619)) ;
    nand02 ix3618 (.Y (nx3617), .A0 (nx314), .A1 (nx5488)) ;
    xnor2 ix3620 (.Y (nx3619), .A0 (nx3621), .A1 (nx3623)) ;
    mux21 ix3622 (.Y (nx3621), .A0 (nx3489), .A1 (nx3495), .S0 (nx3491)) ;
    xnor2 ix3624 (.Y (nx3623), .A0 (nx3625), .A1 (nx3627)) ;
    nand02 ix3626 (.Y (nx3625), .A0 (nx5484), .A1 (nx290)) ;
    xnor2 ix3628 (.Y (nx3627), .A0 (nx3629), .A1 (nx3631)) ;
    mux21 ix3630 (.Y (nx3629), .A0 (nx3497), .A1 (nx3503), .S0 (nx3499)) ;
    xnor2 ix3632 (.Y (nx3631), .A0 (nx3633), .A1 (nx3635)) ;
    nand02 ix3634 (.Y (nx3633), .A0 (nx5480), .A1 (nx266)) ;
    xnor2 ix3636 (.Y (nx3635), .A0 (nx3637), .A1 (nx3639)) ;
    mux21 ix3638 (.Y (nx3637), .A0 (nx3505), .A1 (nx3511), .S0 (nx3507)) ;
    xnor2 ix3640 (.Y (nx3639), .A0 (nx3641), .A1 (nx3643)) ;
    nand02 ix3642 (.Y (nx3641), .A0 (nx5476), .A1 (nx242)) ;
    xnor2 ix3644 (.Y (nx3643), .A0 (nx3645), .A1 (nx3647)) ;
    mux21 ix3646 (.Y (nx3645), .A0 (nx3513), .A1 (nx3519), .S0 (nx3515)) ;
    xnor2 ix3648 (.Y (nx3647), .A0 (nx3649), .A1 (nx3651)) ;
    nand02 ix3650 (.Y (nx3649), .A0 (nx5472), .A1 (nx218)) ;
    xnor2 ix3652 (.Y (nx3651), .A0 (nx3653), .A1 (nx3655)) ;
    mux21 ix3654 (.Y (nx3653), .A0 (nx3521), .A1 (nx3527), .S0 (nx3523)) ;
    xnor2 ix3656 (.Y (nx3655), .A0 (nx3657), .A1 (nx3659)) ;
    nand02 ix3658 (.Y (nx3657), .A0 (nx5468), .A1 (nx194)) ;
    xnor2 ix3660 (.Y (nx3659), .A0 (nx3661), .A1 (nx3663)) ;
    mux21 ix3662 (.Y (nx3661), .A0 (nx3529), .A1 (nx3535), .S0 (nx3531)) ;
    xnor2 ix3664 (.Y (nx3663), .A0 (nx3665), .A1 (nx3667)) ;
    nand02 ix3666 (.Y (nx3665), .A0 (nx5456), .A1 (nx170)) ;
    nand02 ix3668 (.Y (nx3667), .A0 (nx5448), .A1 (nx146)) ;
    mux21 ix147 (.Y (nx146), .A0 (C[13]), .A1 (lfsr_C_13), .S0 (test_mode)) ;
    nor03 ix3131 (.Y (nx3130), .A0 (nx3571), .A1 (nx5536), .A2 (nx3673)) ;
    nor02ii ix4411 (.Y (mac_output[14]), .A0 (RST), .A1 (nx4406)) ;
    nor02 ix4407 (.Y (nx4406), .A0 (RST), .A1 (nx3681)) ;
    xnor2 ix3682 (.Y (nx3681), .A0 (nx3683), .A1 (nx3687)) ;
    xnor2 ix3684 (.Y (nx3683), .A0 (mac_unit_tempP_14), .A1 (nx3980)) ;
    dffr mac_unit_MR_reg_Q_14 (.Q (mac_unit_tempP_14), .QB (\$dummy [45]), .D (
         nx3968), .CLK (CLK), .R (RST)) ;
    aoi22 ix3688 (.Y (nx3687), .A0 (nx3956), .A1 (mac_unit_tempP_13), .B0 (
          nx1915), .B1 (nx3942)) ;
    aoi21 ix3981 (.Y (nx3980), .A0 (nx3697), .A1 (nx3701), .B0 (nx3352)) ;
    mux21 ix3199 (.Y (nx3198), .A0 (B[14]), .A1 (lfsr_C_1), .S0 (test_mode)) ;
    xnor2 ix3702 (.Y (nx3701), .A0 (nx3130), .A1 (nx3120)) ;
    xnor2 ix3121 (.Y (nx3120), .A0 (nx3705), .A1 (nx3116)) ;
    xnor2 ix3117 (.Y (nx3116), .A0 (nx2912), .A1 (nx3709)) ;
    mux21 ix2913 (.Y (nx2912), .A0 (nx2894), .A1 (nx2908), .S0 (nx2898)) ;
    xnor2 ix3710 (.Y (nx3709), .A0 (nx3711), .A1 (nx3713)) ;
    nand02 ix3712 (.Y (nx3711), .A0 (nx410), .A1 (nx5508)) ;
    xnor2 ix3714 (.Y (nx3713), .A0 (nx3715), .A1 (nx3719)) ;
    mux21 ix3716 (.Y (nx3715), .A0 (nx3717), .A1 (nx3585), .S0 (nx3581)) ;
    xnor2 ix3720 (.Y (nx3719), .A0 (nx3721), .A1 (nx3723)) ;
    nand02 ix3722 (.Y (nx3721), .A0 (nx386), .A1 (nx5504)) ;
    xnor2 ix3724 (.Y (nx3723), .A0 (nx3725), .A1 (nx3727)) ;
    mux21 ix3726 (.Y (nx3725), .A0 (nx3587), .A1 (nx3595), .S0 (nx3591)) ;
    xnor2 ix3728 (.Y (nx3727), .A0 (nx3729), .A1 (nx3731)) ;
    nand02 ix3730 (.Y (nx3729), .A0 (nx362), .A1 (nx5500)) ;
    xnor2 ix3732 (.Y (nx3731), .A0 (nx3733), .A1 (nx3735)) ;
    mux21 ix3734 (.Y (nx3733), .A0 (nx3597), .A1 (nx3603), .S0 (nx3599)) ;
    xnor2 ix3736 (.Y (nx3735), .A0 (nx3737), .A1 (nx3739)) ;
    nand02 ix3738 (.Y (nx3737), .A0 (nx338), .A1 (nx5496)) ;
    xnor2 ix3740 (.Y (nx3739), .A0 (nx3741), .A1 (nx3743)) ;
    mux21 ix3742 (.Y (nx3741), .A0 (nx3605), .A1 (nx3611), .S0 (nx3607)) ;
    xnor2 ix3744 (.Y (nx3743), .A0 (nx3745), .A1 (nx3747)) ;
    nand02 ix3746 (.Y (nx3745), .A0 (nx314), .A1 (nx5492)) ;
    xnor2 ix3748 (.Y (nx3747), .A0 (nx3749), .A1 (nx3751)) ;
    mux21 ix3750 (.Y (nx3749), .A0 (nx3613), .A1 (nx3619), .S0 (nx3615)) ;
    xnor2 ix3752 (.Y (nx3751), .A0 (nx3753), .A1 (nx3755)) ;
    nand02 ix3754 (.Y (nx3753), .A0 (nx5488), .A1 (nx290)) ;
    xnor2 ix3756 (.Y (nx3755), .A0 (nx3757), .A1 (nx3759)) ;
    mux21 ix3758 (.Y (nx3757), .A0 (nx3621), .A1 (nx3627), .S0 (nx3623)) ;
    xnor2 ix3760 (.Y (nx3759), .A0 (nx3761), .A1 (nx3763)) ;
    nand02 ix3762 (.Y (nx3761), .A0 (nx5484), .A1 (nx266)) ;
    xnor2 ix3764 (.Y (nx3763), .A0 (nx3765), .A1 (nx3767)) ;
    mux21 ix3766 (.Y (nx3765), .A0 (nx3629), .A1 (nx3635), .S0 (nx3631)) ;
    xnor2 ix3768 (.Y (nx3767), .A0 (nx3769), .A1 (nx3771)) ;
    nand02 ix3770 (.Y (nx3769), .A0 (nx5480), .A1 (nx242)) ;
    xnor2 ix3772 (.Y (nx3771), .A0 (nx3773), .A1 (nx3775)) ;
    mux21 ix3774 (.Y (nx3773), .A0 (nx3637), .A1 (nx3643), .S0 (nx3639)) ;
    xnor2 ix3776 (.Y (nx3775), .A0 (nx3777), .A1 (nx3779)) ;
    nand02 ix3778 (.Y (nx3777), .A0 (nx5476), .A1 (nx218)) ;
    xnor2 ix3780 (.Y (nx3779), .A0 (nx3781), .A1 (nx3783)) ;
    mux21 ix3782 (.Y (nx3781), .A0 (nx3645), .A1 (nx3651), .S0 (nx3647)) ;
    xnor2 ix3784 (.Y (nx3783), .A0 (nx3785), .A1 (nx3787)) ;
    nand02 ix3786 (.Y (nx3785), .A0 (nx5472), .A1 (nx194)) ;
    xnor2 ix3788 (.Y (nx3787), .A0 (nx3789), .A1 (nx3791)) ;
    mux21 ix3790 (.Y (nx3789), .A0 (nx3653), .A1 (nx3659), .S0 (nx3655)) ;
    xnor2 ix3792 (.Y (nx3791), .A0 (nx3793), .A1 (nx3795)) ;
    nand02 ix3794 (.Y (nx3793), .A0 (nx5468), .A1 (nx170)) ;
    xnor2 ix3796 (.Y (nx3795), .A0 (nx3797), .A1 (nx3799)) ;
    mux21 ix3798 (.Y (nx3797), .A0 (nx3661), .A1 (nx3667), .S0 (nx3663)) ;
    xnor2 ix3800 (.Y (nx3799), .A0 (nx3801), .A1 (nx3803)) ;
    nand02 ix3802 (.Y (nx3801), .A0 (nx5456), .A1 (nx146)) ;
    nand02 ix3804 (.Y (nx3803), .A0 (nx5450), .A1 (nx122)) ;
    mux21 ix123 (.Y (nx122), .A0 (C[14]), .A1 (lfsr_C_14), .S0 (test_mode)) ;
    nor03 ix3353 (.Y (nx3352), .A0 (nx3701), .A1 (nx5536), .A2 (nx3807)) ;
    nor02ii ix4419 (.Y (mac_output[15]), .A0 (RST), .A1 (nx4414)) ;
    nor02 ix4415 (.Y (nx4414), .A0 (RST), .A1 (nx3815)) ;
    xnor2 ix3816 (.Y (nx3815), .A0 (nx3817), .A1 (nx3823)) ;
    xnor2 ix3818 (.Y (nx3817), .A0 (mac_unit_tempP_15), .A1 (nx4004)) ;
    dffr mac_unit_MR_reg_Q_15 (.Q (mac_unit_tempP_15), .QB (\$dummy [46]), .D (
         nx3992), .CLK (CLK), .R (RST)) ;
    aoi22 ix3824 (.Y (nx3823), .A0 (nx3980), .A1 (mac_unit_tempP_14), .B0 (
          nx1913), .B1 (nx3966)) ;
    aoi21 ix4005 (.Y (nx4004), .A0 (nx3833), .A1 (nx3837), .B0 (nx3574)) ;
    mux21 ix3421 (.Y (nx3420), .A0 (B[15]), .A1 (lfsr_B_15), .S0 (test_mode)) ;
    xnor2 ix3838 (.Y (nx3837), .A0 (nx3352), .A1 (nx3342)) ;
    xnor2 ix3343 (.Y (nx3342), .A0 (nx3841), .A1 (nx3338)) ;
    xnor2 ix3339 (.Y (nx3338), .A0 (nx3134), .A1 (nx3847)) ;
    mux21 ix3135 (.Y (nx3134), .A0 (nx3116), .A1 (nx3130), .S0 (nx3120)) ;
    xnor2 ix3848 (.Y (nx3847), .A0 (nx3849), .A1 (nx3851)) ;
    nand02 ix3850 (.Y (nx3849), .A0 (nx410), .A1 (nx5512)) ;
    xnor2 ix3852 (.Y (nx3851), .A0 (nx3853), .A1 (nx3857)) ;
    mux21 ix3854 (.Y (nx3853), .A0 (nx3855), .A1 (nx3713), .S0 (nx3709)) ;
    xnor2 ix3858 (.Y (nx3857), .A0 (nx3859), .A1 (nx3861)) ;
    nand02 ix3860 (.Y (nx3859), .A0 (nx386), .A1 (nx5508)) ;
    xnor2 ix3862 (.Y (nx3861), .A0 (nx3863), .A1 (nx3865)) ;
    mux21 ix3864 (.Y (nx3863), .A0 (nx3715), .A1 (nx3723), .S0 (nx3719)) ;
    xnor2 ix3866 (.Y (nx3865), .A0 (nx3867), .A1 (nx3869)) ;
    nand02 ix3868 (.Y (nx3867), .A0 (nx362), .A1 (nx5504)) ;
    xnor2 ix3870 (.Y (nx3869), .A0 (nx3871), .A1 (nx3873)) ;
    mux21 ix3872 (.Y (nx3871), .A0 (nx3725), .A1 (nx3731), .S0 (nx3727)) ;
    xnor2 ix3874 (.Y (nx3873), .A0 (nx3875), .A1 (nx3877)) ;
    nand02 ix3876 (.Y (nx3875), .A0 (nx338), .A1 (nx5500)) ;
    xnor2 ix3878 (.Y (nx3877), .A0 (nx3879), .A1 (nx3881)) ;
    mux21 ix3880 (.Y (nx3879), .A0 (nx3733), .A1 (nx3739), .S0 (nx3735)) ;
    xnor2 ix3882 (.Y (nx3881), .A0 (nx3883), .A1 (nx3885)) ;
    nand02 ix3884 (.Y (nx3883), .A0 (nx314), .A1 (nx5496)) ;
    xnor2 ix3886 (.Y (nx3885), .A0 (nx3887), .A1 (nx3889)) ;
    mux21 ix3888 (.Y (nx3887), .A0 (nx3741), .A1 (nx3747), .S0 (nx3743)) ;
    xnor2 ix3890 (.Y (nx3889), .A0 (nx3891), .A1 (nx3893)) ;
    nand02 ix3892 (.Y (nx3891), .A0 (nx290), .A1 (nx5492)) ;
    xnor2 ix3894 (.Y (nx3893), .A0 (nx3895), .A1 (nx3897)) ;
    mux21 ix3896 (.Y (nx3895), .A0 (nx3749), .A1 (nx3755), .S0 (nx3751)) ;
    xnor2 ix3898 (.Y (nx3897), .A0 (nx3899), .A1 (nx3901)) ;
    nand02 ix3900 (.Y (nx3899), .A0 (nx5488), .A1 (nx266)) ;
    xnor2 ix3902 (.Y (nx3901), .A0 (nx3903), .A1 (nx3905)) ;
    mux21 ix3904 (.Y (nx3903), .A0 (nx3757), .A1 (nx3763), .S0 (nx3759)) ;
    xnor2 ix3906 (.Y (nx3905), .A0 (nx3907), .A1 (nx3909)) ;
    nand02 ix3908 (.Y (nx3907), .A0 (nx5484), .A1 (nx242)) ;
    xnor2 ix3910 (.Y (nx3909), .A0 (nx3911), .A1 (nx3913)) ;
    mux21 ix3912 (.Y (nx3911), .A0 (nx3765), .A1 (nx3771), .S0 (nx3767)) ;
    xnor2 ix3914 (.Y (nx3913), .A0 (nx3915), .A1 (nx3917)) ;
    nand02 ix3916 (.Y (nx3915), .A0 (nx5480), .A1 (nx218)) ;
    xnor2 ix3918 (.Y (nx3917), .A0 (nx3919), .A1 (nx3921)) ;
    mux21 ix3920 (.Y (nx3919), .A0 (nx3773), .A1 (nx3779), .S0 (nx3775)) ;
    xnor2 ix3922 (.Y (nx3921), .A0 (nx3923), .A1 (nx3925)) ;
    nand02 ix3924 (.Y (nx3923), .A0 (nx5476), .A1 (nx194)) ;
    xnor2 ix3926 (.Y (nx3925), .A0 (nx3927), .A1 (nx3929)) ;
    mux21 ix3928 (.Y (nx3927), .A0 (nx3781), .A1 (nx3787), .S0 (nx3783)) ;
    xnor2 ix3930 (.Y (nx3929), .A0 (nx3931), .A1 (nx3933)) ;
    nand02 ix3932 (.Y (nx3931), .A0 (nx5472), .A1 (nx170)) ;
    xnor2 ix3934 (.Y (nx3933), .A0 (nx3935), .A1 (nx3937)) ;
    mux21 ix3936 (.Y (nx3935), .A0 (nx3789), .A1 (nx3795), .S0 (nx3791)) ;
    xnor2 ix3938 (.Y (nx3937), .A0 (nx3939), .A1 (nx3941)) ;
    nand02 ix3940 (.Y (nx3939), .A0 (nx5468), .A1 (nx146)) ;
    xnor2 ix3942 (.Y (nx3941), .A0 (nx3943), .A1 (nx3945)) ;
    mux21 ix3944 (.Y (nx3943), .A0 (nx3797), .A1 (nx3803), .S0 (nx3799)) ;
    xnor2 ix3946 (.Y (nx3945), .A0 (nx3947), .A1 (nx3949)) ;
    nand02 ix3948 (.Y (nx3947), .A0 (nx5456), .A1 (nx122)) ;
    mux21 ix99 (.Y (nx98), .A0 (C[15]), .A1 (lfsr_C_15), .S0 (test_mode)) ;
    nor03 ix3575 (.Y (nx3574), .A0 (nx3837), .A1 (nx5536), .A2 (nx3955)) ;
    nor02ii ix4427 (.Y (mac_output[16]), .A0 (RST), .A1 (nx4422)) ;
    nor02 ix4423 (.Y (nx4422), .A0 (RST), .A1 (nx3963)) ;
    xnor2 ix3964 (.Y (nx3963), .A0 (nx3965), .A1 (nx3971)) ;
    xnor2 ix3966 (.Y (nx3965), .A0 (mac_unit_tempP_16), .A1 (nx4022)) ;
    dffr mac_unit_MR_reg_Q_16 (.Q (mac_unit_tempP_16), .QB (\$dummy [47]), .D (
         nx4016), .CLK (CLK), .R (RST)) ;
    aoi22 ix3972 (.Y (nx3971), .A0 (nx4004), .A1 (mac_unit_tempP_15), .B0 (
          nx1912), .B1 (nx3990)) ;
    xnor2 ix4023 (.Y (nx4022), .A0 (nx3574), .A1 (nx3979)) ;
    xnor2 ix3980 (.Y (nx3979), .A0 (nx3981), .A1 (nx3983)) ;
    xnor2 ix3984 (.Y (nx3983), .A0 (nx3356), .A1 (nx3332)) ;
    mux21 ix3357 (.Y (nx3356), .A0 (nx3338), .A1 (nx3352), .S0 (nx3342)) ;
    xnor2 ix3333 (.Y (nx3332), .A0 (nx3989), .A1 (nx3328)) ;
    nand02 ix3990 (.Y (nx3989), .A0 (nx410), .A1 (nx5516)) ;
    xnor2 ix3329 (.Y (nx3328), .A0 (nx3993), .A1 (nx3100)) ;
    mux21 ix3994 (.Y (nx3993), .A0 (nx3995), .A1 (nx3851), .S0 (nx3847)) ;
    xnor2 ix3101 (.Y (nx3100), .A0 (nx3999), .A1 (nx3096)) ;
    nand02 ix4000 (.Y (nx3999), .A0 (nx386), .A1 (nx5512)) ;
    xnor2 ix3097 (.Y (nx3096), .A0 (nx4003), .A1 (nx2868)) ;
    mux21 ix4004 (.Y (nx4003), .A0 (nx3853), .A1 (nx3861), .S0 (nx3857)) ;
    xnor2 ix2869 (.Y (nx2868), .A0 (nx4007), .A1 (nx2864)) ;
    nand02 ix4008 (.Y (nx4007), .A0 (nx362), .A1 (nx5508)) ;
    xnor2 ix2865 (.Y (nx2864), .A0 (nx4011), .A1 (nx2636)) ;
    mux21 ix4012 (.Y (nx4011), .A0 (nx3863), .A1 (nx3869), .S0 (nx3865)) ;
    xnor2 ix2637 (.Y (nx2636), .A0 (nx4015), .A1 (nx2632)) ;
    nand02 ix4016 (.Y (nx4015), .A0 (nx338), .A1 (nx5504)) ;
    xnor2 ix2633 (.Y (nx2632), .A0 (nx4019), .A1 (nx2404)) ;
    mux21 ix4020 (.Y (nx4019), .A0 (nx3871), .A1 (nx3877), .S0 (nx3873)) ;
    xnor2 ix2405 (.Y (nx2404), .A0 (nx4023), .A1 (nx2400)) ;
    nand02 ix4024 (.Y (nx4023), .A0 (nx314), .A1 (nx5500)) ;
    xnor2 ix2401 (.Y (nx2400), .A0 (nx4027), .A1 (nx2172)) ;
    mux21 ix4028 (.Y (nx4027), .A0 (nx3879), .A1 (nx3885), .S0 (nx3881)) ;
    xnor2 ix2173 (.Y (nx2172), .A0 (nx4031), .A1 (nx2168)) ;
    nand02 ix4032 (.Y (nx4031), .A0 (nx290), .A1 (nx5496)) ;
    xnor2 ix2169 (.Y (nx2168), .A0 (nx4035), .A1 (nx1940)) ;
    mux21 ix4036 (.Y (nx4035), .A0 (nx3887), .A1 (nx3893), .S0 (nx3889)) ;
    xnor2 ix1941 (.Y (nx1940), .A0 (nx4038), .A1 (nx1936)) ;
    nand02 ix4039 (.Y (nx4038), .A0 (nx5492), .A1 (nx266)) ;
    xnor2 ix1937 (.Y (nx1936), .A0 (nx4041), .A1 (nx1708)) ;
    mux21 ix4042 (.Y (nx4041), .A0 (nx3895), .A1 (nx3901), .S0 (nx3897)) ;
    xnor2 ix1709 (.Y (nx1708), .A0 (nx4045), .A1 (nx1704)) ;
    nand02 ix4046 (.Y (nx4045), .A0 (nx5488), .A1 (nx242)) ;
    xnor2 ix1705 (.Y (nx1704), .A0 (nx4049), .A1 (nx1476)) ;
    mux21 ix4050 (.Y (nx4049), .A0 (nx3903), .A1 (nx3909), .S0 (nx3905)) ;
    xnor2 ix1477 (.Y (nx1476), .A0 (nx4053), .A1 (nx1472)) ;
    nand02 ix4054 (.Y (nx4053), .A0 (nx5484), .A1 (nx218)) ;
    xnor2 ix1473 (.Y (nx1472), .A0 (nx4056), .A1 (nx1244)) ;
    mux21 ix4057 (.Y (nx4056), .A0 (nx3911), .A1 (nx3917), .S0 (nx3913)) ;
    xnor2 ix1245 (.Y (nx1244), .A0 (nx4059), .A1 (nx1240)) ;
    nand02 ix4060 (.Y (nx4059), .A0 (nx5480), .A1 (nx194)) ;
    xnor2 ix1241 (.Y (nx1240), .A0 (nx4063), .A1 (nx1012)) ;
    mux21 ix4064 (.Y (nx4063), .A0 (nx3919), .A1 (nx3925), .S0 (nx3921)) ;
    xnor2 ix1013 (.Y (nx1012), .A0 (nx4067), .A1 (nx1008)) ;
    nand02 ix4068 (.Y (nx4067), .A0 (nx5476), .A1 (nx170)) ;
    xnor2 ix1009 (.Y (nx1008), .A0 (nx4071), .A1 (nx780)) ;
    mux21 ix4072 (.Y (nx4071), .A0 (nx3927), .A1 (nx3933), .S0 (nx3929)) ;
    xnor2 ix781 (.Y (nx780), .A0 (nx4074), .A1 (nx776)) ;
    nand02 ix4075 (.Y (nx4074), .A0 (nx5472), .A1 (nx146)) ;
    xnor2 ix777 (.Y (nx776), .A0 (nx4077), .A1 (nx548)) ;
    mux21 ix4078 (.Y (nx4077), .A0 (nx3935), .A1 (nx3941), .S0 (nx3937)) ;
    xnor2 ix549 (.Y (nx548), .A0 (nx4081), .A1 (nx544)) ;
    nand02 ix4082 (.Y (nx4081), .A0 (nx5468), .A1 (nx122)) ;
    aoi21 ix545 (.Y (nx544), .A0 (nx4085), .A1 (nx4087), .B0 (nx520)) ;
    mux21 ix4088 (.Y (nx4087), .A0 (nx3943), .A1 (nx3949), .S0 (nx3945)) ;
    nor03 ix521 (.Y (nx520), .A0 (nx4087), .A1 (nx2583), .A2 (nx5550)) ;
    nor02 ix4435 (.Y (mac_output[17]), .A0 (RST), .A1 (nx4095)) ;
    nand02 ix4096 (.Y (nx4095), .A0 (nx2523), .A1 (nx4034)) ;
    xnor2 ix4035 (.Y (nx4034), .A0 (nx1909), .A1 (nx4239)) ;
    xnor2 ix4043 (.Y (nx1909), .A0 (mac_unit_tempP_17), .A1 (nx4105)) ;
    dffr mac_unit_MR_reg_Q_17 (.Q (mac_unit_tempP_17), .QB (\$dummy [48]), .D (
         nx4034), .CLK (CLK), .R (RST)) ;
    xnor2 ix4106 (.Y (nx4105), .A0 (nx4107), .A1 (nx4111)) ;
    mux21 ix4108 (.Y (nx4107), .A0 (nx4109), .A1 (nx3983), .S0 (nx3979)) ;
    xnor2 ix4112 (.Y (nx4111), .A0 (nx4113), .A1 (nx4115)) ;
    nand02 ix4114 (.Y (nx4113), .A0 (nx410), .A1 (nx5520)) ;
    xnor2 ix4116 (.Y (nx4115), .A0 (nx3360), .A1 (nx3322)) ;
    mux21 ix3361 (.Y (nx3360), .A0 (nx3328), .A1 (nx3356), .S0 (nx3332)) ;
    xnor2 ix3323 (.Y (nx3322), .A0 (nx4121), .A1 (nx3318)) ;
    nand02 ix4122 (.Y (nx4121), .A0 (nx386), .A1 (nx5516)) ;
    xnor2 ix3319 (.Y (nx3318), .A0 (nx4125), .A1 (nx3090)) ;
    mux21 ix4126 (.Y (nx4125), .A0 (nx4127), .A1 (nx3993), .S0 (nx3100)) ;
    xnor2 ix3091 (.Y (nx3090), .A0 (nx4131), .A1 (nx3086)) ;
    nand02 ix4132 (.Y (nx4131), .A0 (nx362), .A1 (nx5512)) ;
    xnor2 ix3087 (.Y (nx3086), .A0 (nx4135), .A1 (nx2858)) ;
    mux21 ix4136 (.Y (nx4135), .A0 (nx4137), .A1 (nx4003), .S0 (nx2868)) ;
    xnor2 ix2859 (.Y (nx2858), .A0 (nx4141), .A1 (nx2854)) ;
    nand02 ix4142 (.Y (nx4141), .A0 (nx338), .A1 (nx5508)) ;
    xnor2 ix2855 (.Y (nx2854), .A0 (nx4145), .A1 (nx2626)) ;
    mux21 ix4146 (.Y (nx4145), .A0 (nx4147), .A1 (nx4011), .S0 (nx2636)) ;
    xnor2 ix2627 (.Y (nx2626), .A0 (nx4151), .A1 (nx2622)) ;
    nand02 ix4152 (.Y (nx4151), .A0 (nx314), .A1 (nx5504)) ;
    xnor2 ix2623 (.Y (nx2622), .A0 (nx4155), .A1 (nx2394)) ;
    mux21 ix4156 (.Y (nx4155), .A0 (nx4157), .A1 (nx4019), .S0 (nx2404)) ;
    xnor2 ix2395 (.Y (nx2394), .A0 (nx4161), .A1 (nx2390)) ;
    nand02 ix4162 (.Y (nx4161), .A0 (nx290), .A1 (nx5500)) ;
    xnor2 ix2391 (.Y (nx2390), .A0 (nx4164), .A1 (nx2162)) ;
    mux21 ix4165 (.Y (nx4164), .A0 (nx4167), .A1 (nx4027), .S0 (nx2172)) ;
    xnor2 ix2163 (.Y (nx2162), .A0 (nx4171), .A1 (nx2158)) ;
    nand02 ix4172 (.Y (nx4171), .A0 (nx266), .A1 (nx5496)) ;
    xnor2 ix2159 (.Y (nx2158), .A0 (nx4175), .A1 (nx1930)) ;
    mux21 ix4176 (.Y (nx4175), .A0 (nx4177), .A1 (nx4035), .S0 (nx1940)) ;
    xnor2 ix1931 (.Y (nx1930), .A0 (nx4181), .A1 (nx1926)) ;
    nand02 ix4182 (.Y (nx4181), .A0 (nx5492), .A1 (nx242)) ;
    xnor2 ix1927 (.Y (nx1926), .A0 (nx4185), .A1 (nx1698)) ;
    mux21 ix4186 (.Y (nx4185), .A0 (nx4187), .A1 (nx4041), .S0 (nx1708)) ;
    xnor2 ix1699 (.Y (nx1698), .A0 (nx4191), .A1 (nx1694)) ;
    nand02 ix4192 (.Y (nx4191), .A0 (nx5488), .A1 (nx218)) ;
    xnor2 ix1695 (.Y (nx1694), .A0 (nx4195), .A1 (nx1466)) ;
    mux21 ix4196 (.Y (nx4195), .A0 (nx4197), .A1 (nx4049), .S0 (nx1476)) ;
    xnor2 ix1467 (.Y (nx1466), .A0 (nx4200), .A1 (nx1462)) ;
    nand02 ix4201 (.Y (nx4200), .A0 (nx5484), .A1 (nx194)) ;
    xnor2 ix1463 (.Y (nx1462), .A0 (nx4203), .A1 (nx1234)) ;
    mux21 ix4204 (.Y (nx4203), .A0 (nx4205), .A1 (nx4056), .S0 (nx1244)) ;
    xnor2 ix1235 (.Y (nx1234), .A0 (nx4209), .A1 (nx1230)) ;
    nand02 ix4210 (.Y (nx4209), .A0 (nx5480), .A1 (nx170)) ;
    xnor2 ix1231 (.Y (nx1230), .A0 (nx4213), .A1 (nx1002)) ;
    mux21 ix4214 (.Y (nx4213), .A0 (nx4215), .A1 (nx4063), .S0 (nx1012)) ;
    xnor2 ix1003 (.Y (nx1002), .A0 (nx4218), .A1 (nx998)) ;
    nand02 ix4219 (.Y (nx4218), .A0 (nx5476), .A1 (nx146)) ;
    xnor2 ix999 (.Y (nx998), .A0 (nx4221), .A1 (nx770)) ;
    mux21 ix4222 (.Y (nx4221), .A0 (nx4223), .A1 (nx4071), .S0 (nx780)) ;
    xnor2 ix771 (.Y (nx770), .A0 (nx4227), .A1 (nx766)) ;
    nand02 ix4228 (.Y (nx4227), .A0 (nx5472), .A1 (nx122)) ;
    xnor2 ix767 (.Y (nx766), .A0 (nx4231), .A1 (nx532)) ;
    mux21 ix4232 (.Y (nx4231), .A0 (nx4233), .A1 (nx4077), .S0 (nx548)) ;
    xnor2 ix533 (.Y (nx532), .A0 (nx4237), .A1 (nx520)) ;
    aoi22 ix4240 (.Y (nx4239), .A0 (nx4022), .A1 (mac_unit_tempP_16), .B0 (
          nx1911), .B1 (nx4014)) ;
    nor02ii ix4443 (.Y (mac_output[18]), .A0 (RST), .A1 (nx4438)) ;
    nor02 ix4439 (.Y (nx4438), .A0 (RST), .A1 (nx4251)) ;
    xnor2 ix4252 (.Y (nx4251), .A0 (nx4253), .A1 (nx4257)) ;
    xnor2 ix4254 (.Y (nx4253), .A0 (mac_unit_tempP_18), .A1 (nx4058)) ;
    dffr mac_unit_MR_reg_Q_18 (.Q (mac_unit_tempP_18), .QB (\$dummy [49]), .D (
         nx4052), .CLK (CLK), .R (RST)) ;
    mux21 ix4258 (.Y (nx4257), .A0 (nx4105), .A1 (nx4239), .S0 (nx1909)) ;
    xnor2 ix4059 (.Y (nx4058), .A0 (nx4261), .A1 (nx3544)) ;
    mux21 ix4262 (.Y (nx4261), .A0 (nx4107), .A1 (nx4115), .S0 (nx4111)) ;
    xnor2 ix3545 (.Y (nx3544), .A0 (nx4265), .A1 (nx3540)) ;
    nand02 ix4266 (.Y (nx4265), .A0 (nx386), .A1 (nx5520)) ;
    xnor2 ix3541 (.Y (nx3540), .A0 (nx3364), .A1 (nx4271)) ;
    mux21 ix3365 (.Y (nx3364), .A0 (nx3318), .A1 (nx3360), .S0 (nx3322)) ;
    xnor2 ix4272 (.Y (nx4271), .A0 (nx4273), .A1 (nx4275)) ;
    nand02 ix4274 (.Y (nx4273), .A0 (nx362), .A1 (nx5516)) ;
    xnor2 ix4276 (.Y (nx4275), .A0 (nx4277), .A1 (nx4281)) ;
    mux21 ix4278 (.Y (nx4277), .A0 (nx4279), .A1 (nx4125), .S0 (nx3090)) ;
    xnor2 ix4282 (.Y (nx4281), .A0 (nx4283), .A1 (nx4285)) ;
    nand02 ix4284 (.Y (nx4283), .A0 (nx338), .A1 (nx5512)) ;
    xnor2 ix4286 (.Y (nx4285), .A0 (nx4287), .A1 (nx4291)) ;
    mux21 ix4288 (.Y (nx4287), .A0 (nx4289), .A1 (nx4135), .S0 (nx2858)) ;
    xnor2 ix4292 (.Y (nx4291), .A0 (nx4293), .A1 (nx4295)) ;
    nand02 ix4294 (.Y (nx4293), .A0 (nx314), .A1 (nx5508)) ;
    xnor2 ix4296 (.Y (nx4295), .A0 (nx4297), .A1 (nx4301)) ;
    mux21 ix4298 (.Y (nx4297), .A0 (nx4299), .A1 (nx4145), .S0 (nx2626)) ;
    xnor2 ix4302 (.Y (nx4301), .A0 (nx4303), .A1 (nx4305)) ;
    nand02 ix4304 (.Y (nx4303), .A0 (nx290), .A1 (nx5504)) ;
    xnor2 ix4306 (.Y (nx4305), .A0 (nx4307), .A1 (nx4311)) ;
    mux21 ix4308 (.Y (nx4307), .A0 (nx4309), .A1 (nx4155), .S0 (nx2394)) ;
    xnor2 ix4312 (.Y (nx4311), .A0 (nx4313), .A1 (nx4315)) ;
    nand02 ix4314 (.Y (nx4313), .A0 (nx266), .A1 (nx5500)) ;
    xnor2 ix4316 (.Y (nx4315), .A0 (nx4317), .A1 (nx4321)) ;
    mux21 ix4318 (.Y (nx4317), .A0 (nx4319), .A1 (nx4164), .S0 (nx2162)) ;
    xnor2 ix4322 (.Y (nx4321), .A0 (nx4323), .A1 (nx4325)) ;
    nand02 ix4324 (.Y (nx4323), .A0 (nx5496), .A1 (nx242)) ;
    xnor2 ix4326 (.Y (nx4325), .A0 (nx4327), .A1 (nx4331)) ;
    mux21 ix4328 (.Y (nx4327), .A0 (nx4329), .A1 (nx4175), .S0 (nx1930)) ;
    xnor2 ix4332 (.Y (nx4331), .A0 (nx4333), .A1 (nx4335)) ;
    nand02 ix4334 (.Y (nx4333), .A0 (nx5492), .A1 (nx218)) ;
    xnor2 ix4336 (.Y (nx4335), .A0 (nx4337), .A1 (nx4341)) ;
    mux21 ix4338 (.Y (nx4337), .A0 (nx4339), .A1 (nx4185), .S0 (nx1698)) ;
    xnor2 ix4342 (.Y (nx4341), .A0 (nx4343), .A1 (nx4345)) ;
    nand02 ix4344 (.Y (nx4343), .A0 (nx5488), .A1 (nx194)) ;
    xnor2 ix4346 (.Y (nx4345), .A0 (nx4347), .A1 (nx4351)) ;
    mux21 ix4348 (.Y (nx4347), .A0 (nx4349), .A1 (nx4195), .S0 (nx1466)) ;
    xnor2 ix4352 (.Y (nx4351), .A0 (nx4353), .A1 (nx4355)) ;
    nand02 ix4354 (.Y (nx4353), .A0 (nx5484), .A1 (nx170)) ;
    xnor2 ix4356 (.Y (nx4355), .A0 (nx4357), .A1 (nx4361)) ;
    mux21 ix4358 (.Y (nx4357), .A0 (nx4359), .A1 (nx4203), .S0 (nx1234)) ;
    xnor2 ix4362 (.Y (nx4361), .A0 (nx4363), .A1 (nx4365)) ;
    nand02 ix4364 (.Y (nx4363), .A0 (nx5480), .A1 (nx146)) ;
    xnor2 ix4366 (.Y (nx4365), .A0 (nx4367), .A1 (nx4371)) ;
    mux21 ix4368 (.Y (nx4367), .A0 (nx4369), .A1 (nx4213), .S0 (nx1002)) ;
    xnor2 ix4372 (.Y (nx4371), .A0 (nx4373), .A1 (nx4375)) ;
    nand02 ix4374 (.Y (nx4373), .A0 (nx5476), .A1 (nx122)) ;
    xnor2 ix4376 (.Y (nx4375), .A0 (nx4377), .A1 (nx4381)) ;
    mux21 ix4378 (.Y (nx4377), .A0 (nx4379), .A1 (nx4221), .S0 (nx770)) ;
    xnor2 ix4382 (.Y (nx4381), .A0 (nx4383), .A1 (nx4385)) ;
    mux21 ix4386 (.Y (nx4385), .A0 (nx4387), .A1 (nx4231), .S0 (nx532)) ;
    nor02 ix4451 (.Y (mac_output[19]), .A0 (RST), .A1 (nx4391)) ;
    nand02 ix4392 (.Y (nx4391), .A0 (nx2523), .A1 (nx4070)) ;
    xnor2 ix4071 (.Y (nx4070), .A0 (nx1905), .A1 (nx4501)) ;
    xnor2 ix4079 (.Y (nx1905), .A0 (mac_unit_tempP_19), .A1 (nx4399)) ;
    dffr mac_unit_MR_reg_Q_19 (.Q (mac_unit_tempP_19), .QB (\$dummy [50]), .D (
         nx4070), .CLK (CLK), .R (RST)) ;
    xnor2 ix4400 (.Y (nx4399), .A0 (nx4401), .A1 (nx4405)) ;
    mux21 ix4402 (.Y (nx4401), .A0 (nx4403), .A1 (nx4261), .S0 (nx3544)) ;
    xnor2 ix4406 (.Y (nx4405), .A0 (nx4407), .A1 (nx4409)) ;
    nand02 ix4408 (.Y (nx4407), .A0 (nx362), .A1 (nx5520)) ;
    xnor2 ix4410 (.Y (nx4409), .A0 (nx4411), .A1 (nx4415)) ;
    mux21 ix4412 (.Y (nx4411), .A0 (nx4413), .A1 (nx4275), .S0 (nx4271)) ;
    xnor2 ix4416 (.Y (nx4415), .A0 (nx4417), .A1 (nx4419)) ;
    nand02 ix4418 (.Y (nx4417), .A0 (nx338), .A1 (nx5516)) ;
    xnor2 ix4420 (.Y (nx4419), .A0 (nx4421), .A1 (nx4423)) ;
    mux21 ix4422 (.Y (nx4421), .A0 (nx4277), .A1 (nx4285), .S0 (nx4281)) ;
    xnor2 ix4424 (.Y (nx4423), .A0 (nx4425), .A1 (nx4427)) ;
    nand02 ix4426 (.Y (nx4425), .A0 (nx314), .A1 (nx5512)) ;
    xnor2 ix4428 (.Y (nx4427), .A0 (nx4429), .A1 (nx4431)) ;
    mux21 ix4430 (.Y (nx4429), .A0 (nx4287), .A1 (nx4295), .S0 (nx4291)) ;
    xnor2 ix4432 (.Y (nx4431), .A0 (nx4433), .A1 (nx4435)) ;
    nand02 ix4434 (.Y (nx4433), .A0 (nx290), .A1 (nx5508)) ;
    xnor2 ix4436 (.Y (nx4435), .A0 (nx4437), .A1 (nx4439)) ;
    mux21 ix4438 (.Y (nx4437), .A0 (nx4297), .A1 (nx4305), .S0 (nx4301)) ;
    xnor2 ix4440 (.Y (nx4439), .A0 (nx4441), .A1 (nx4443)) ;
    nand02 ix4442 (.Y (nx4441), .A0 (nx266), .A1 (nx5504)) ;
    xnor2 ix4444 (.Y (nx4443), .A0 (nx4445), .A1 (nx4447)) ;
    mux21 ix4446 (.Y (nx4445), .A0 (nx4307), .A1 (nx4315), .S0 (nx4311)) ;
    xnor2 ix4448 (.Y (nx4447), .A0 (nx4449), .A1 (nx4451)) ;
    nand02 ix4450 (.Y (nx4449), .A0 (nx242), .A1 (nx5500)) ;
    xnor2 ix4452 (.Y (nx4451), .A0 (nx4453), .A1 (nx4455)) ;
    mux21 ix4454 (.Y (nx4453), .A0 (nx4317), .A1 (nx4325), .S0 (nx4321)) ;
    xnor2 ix4456 (.Y (nx4455), .A0 (nx4457), .A1 (nx4459)) ;
    nand02 ix4458 (.Y (nx4457), .A0 (nx5496), .A1 (nx218)) ;
    xnor2 ix4460 (.Y (nx4459), .A0 (nx4461), .A1 (nx4463)) ;
    mux21 ix4462 (.Y (nx4461), .A0 (nx4327), .A1 (nx4335), .S0 (nx4331)) ;
    xnor2 ix4464 (.Y (nx4463), .A0 (nx4465), .A1 (nx4467)) ;
    nand02 ix4466 (.Y (nx4465), .A0 (nx5492), .A1 (nx194)) ;
    xnor2 ix4468 (.Y (nx4467), .A0 (nx4469), .A1 (nx4471)) ;
    mux21 ix4470 (.Y (nx4469), .A0 (nx4337), .A1 (nx4345), .S0 (nx4341)) ;
    xnor2 ix4472 (.Y (nx4471), .A0 (nx4473), .A1 (nx4475)) ;
    nand02 ix4474 (.Y (nx4473), .A0 (nx5488), .A1 (nx170)) ;
    xnor2 ix4476 (.Y (nx4475), .A0 (nx4477), .A1 (nx4479)) ;
    mux21 ix4478 (.Y (nx4477), .A0 (nx4347), .A1 (nx4355), .S0 (nx4351)) ;
    xnor2 ix4480 (.Y (nx4479), .A0 (nx4481), .A1 (nx4483)) ;
    nand02 ix4482 (.Y (nx4481), .A0 (nx5484), .A1 (nx146)) ;
    xnor2 ix4484 (.Y (nx4483), .A0 (nx4485), .A1 (nx4487)) ;
    mux21 ix4486 (.Y (nx4485), .A0 (nx4357), .A1 (nx4365), .S0 (nx4361)) ;
    xnor2 ix4488 (.Y (nx4487), .A0 (nx4489), .A1 (nx4491)) ;
    nand02 ix4490 (.Y (nx4489), .A0 (nx5480), .A1 (nx122)) ;
    xnor2 ix4492 (.Y (nx4491), .A0 (nx4493), .A1 (nx4495)) ;
    mux21 ix4494 (.Y (nx4493), .A0 (nx4367), .A1 (nx4375), .S0 (nx4371)) ;
    xnor2 ix4496 (.Y (nx4495), .A0 (nx4497), .A1 (nx4499)) ;
    mux21 ix4500 (.Y (nx4499), .A0 (nx4377), .A1 (nx4385), .S0 (nx4381)) ;
    aoi22 ix4502 (.Y (nx4501), .A0 (nx4058), .A1 (mac_unit_tempP_18), .B0 (
          nx1907), .B1 (nx4050)) ;
    nor02 ix4459 (.Y (mac_output[20]), .A0 (RST), .A1 (nx4511)) ;
    nand02 ix4512 (.Y (nx4511), .A0 (nx2523), .A1 (nx4088)) ;
    xnor2 ix4089 (.Y (nx4088), .A0 (nx1903), .A1 (nx4609)) ;
    xnor2 ix4097 (.Y (nx1903), .A0 (mac_unit_tempP_20), .A1 (nx4519)) ;
    dffr mac_unit_MR_reg_Q_20 (.Q (mac_unit_tempP_20), .QB (\$dummy [51]), .D (
         nx4088), .CLK (CLK), .R (RST)) ;
    xnor2 ix4520 (.Y (nx4519), .A0 (nx4521), .A1 (nx4523)) ;
    mux21 ix4522 (.Y (nx4521), .A0 (nx4401), .A1 (nx4409), .S0 (nx4405)) ;
    xnor2 ix4524 (.Y (nx4523), .A0 (nx4525), .A1 (nx4527)) ;
    nand02 ix4526 (.Y (nx4525), .A0 (nx338), .A1 (nx5520)) ;
    xnor2 ix4528 (.Y (nx4527), .A0 (nx4529), .A1 (nx4531)) ;
    mux21 ix4530 (.Y (nx4529), .A0 (nx4411), .A1 (nx4419), .S0 (nx4415)) ;
    xnor2 ix4532 (.Y (nx4531), .A0 (nx4533), .A1 (nx4535)) ;
    nand02 ix4534 (.Y (nx4533), .A0 (nx314), .A1 (nx5516)) ;
    xnor2 ix4536 (.Y (nx4535), .A0 (nx4537), .A1 (nx4539)) ;
    mux21 ix4538 (.Y (nx4537), .A0 (nx4421), .A1 (nx4427), .S0 (nx4423)) ;
    xnor2 ix4540 (.Y (nx4539), .A0 (nx4541), .A1 (nx4543)) ;
    nand02 ix4542 (.Y (nx4541), .A0 (nx290), .A1 (nx5512)) ;
    xnor2 ix4544 (.Y (nx4543), .A0 (nx4545), .A1 (nx4547)) ;
    mux21 ix4546 (.Y (nx4545), .A0 (nx4429), .A1 (nx4435), .S0 (nx4431)) ;
    xnor2 ix4548 (.Y (nx4547), .A0 (nx4549), .A1 (nx4551)) ;
    nand02 ix4550 (.Y (nx4549), .A0 (nx266), .A1 (nx5508)) ;
    xnor2 ix4552 (.Y (nx4551), .A0 (nx4553), .A1 (nx4555)) ;
    mux21 ix4554 (.Y (nx4553), .A0 (nx4437), .A1 (nx4443), .S0 (nx4439)) ;
    xnor2 ix4556 (.Y (nx4555), .A0 (nx4557), .A1 (nx4559)) ;
    nand02 ix4558 (.Y (nx4557), .A0 (nx242), .A1 (nx5504)) ;
    xnor2 ix4560 (.Y (nx4559), .A0 (nx4561), .A1 (nx4563)) ;
    mux21 ix4562 (.Y (nx4561), .A0 (nx4445), .A1 (nx4451), .S0 (nx4447)) ;
    xnor2 ix4564 (.Y (nx4563), .A0 (nx4565), .A1 (nx4567)) ;
    nand02 ix4566 (.Y (nx4565), .A0 (nx5500), .A1 (nx218)) ;
    xnor2 ix4568 (.Y (nx4567), .A0 (nx4569), .A1 (nx4571)) ;
    mux21 ix4570 (.Y (nx4569), .A0 (nx4453), .A1 (nx4459), .S0 (nx4455)) ;
    xnor2 ix4572 (.Y (nx4571), .A0 (nx4573), .A1 (nx4575)) ;
    nand02 ix4574 (.Y (nx4573), .A0 (nx5496), .A1 (nx194)) ;
    xnor2 ix4576 (.Y (nx4575), .A0 (nx4577), .A1 (nx4579)) ;
    mux21 ix4578 (.Y (nx4577), .A0 (nx4461), .A1 (nx4467), .S0 (nx4463)) ;
    xnor2 ix4580 (.Y (nx4579), .A0 (nx4581), .A1 (nx4583)) ;
    nand02 ix4582 (.Y (nx4581), .A0 (nx5492), .A1 (nx170)) ;
    xnor2 ix4584 (.Y (nx4583), .A0 (nx4585), .A1 (nx4587)) ;
    mux21 ix4586 (.Y (nx4585), .A0 (nx4469), .A1 (nx4475), .S0 (nx4471)) ;
    xnor2 ix4588 (.Y (nx4587), .A0 (nx4589), .A1 (nx4591)) ;
    nand02 ix4590 (.Y (nx4589), .A0 (nx5488), .A1 (nx146)) ;
    xnor2 ix4592 (.Y (nx4591), .A0 (nx4593), .A1 (nx4595)) ;
    mux21 ix4594 (.Y (nx4593), .A0 (nx4477), .A1 (nx4483), .S0 (nx4479)) ;
    xnor2 ix4596 (.Y (nx4595), .A0 (nx4597), .A1 (nx4599)) ;
    nand02 ix4598 (.Y (nx4597), .A0 (nx5484), .A1 (nx122)) ;
    xnor2 ix4600 (.Y (nx4599), .A0 (nx4601), .A1 (nx4603)) ;
    mux21 ix4602 (.Y (nx4601), .A0 (nx4485), .A1 (nx4491), .S0 (nx4487)) ;
    xnor2 ix4604 (.Y (nx4603), .A0 (nx4605), .A1 (nx4607)) ;
    mux21 ix4608 (.Y (nx4607), .A0 (nx4493), .A1 (nx4499), .S0 (nx4495)) ;
    mux21 ix4610 (.Y (nx4609), .A0 (nx4399), .A1 (nx4501), .S0 (nx1905)) ;
    nor02 ix4467 (.Y (mac_output[21]), .A0 (RST), .A1 (nx4613)) ;
    nand02 ix4614 (.Y (nx4613), .A0 (nx2523), .A1 (nx4106)) ;
    xnor2 ix4107 (.Y (nx4106), .A0 (nx1902), .A1 (nx4703)) ;
    xnor2 ix4115 (.Y (nx1902), .A0 (mac_unit_tempP_21), .A1 (nx4620)) ;
    dffr mac_unit_MR_reg_Q_21 (.Q (mac_unit_tempP_21), .QB (\$dummy [52]), .D (
         nx4106), .CLK (CLK), .R (RST)) ;
    xnor2 ix4621 (.Y (nx4620), .A0 (nx4623), .A1 (nx4625)) ;
    mux21 ix4624 (.Y (nx4623), .A0 (nx4521), .A1 (nx4527), .S0 (nx4523)) ;
    xnor2 ix4626 (.Y (nx4625), .A0 (nx4627), .A1 (nx4629)) ;
    nand02 ix4628 (.Y (nx4627), .A0 (nx314), .A1 (nx5520)) ;
    xnor2 ix4630 (.Y (nx4629), .A0 (nx4631), .A1 (nx4633)) ;
    mux21 ix4632 (.Y (nx4631), .A0 (nx4529), .A1 (nx4535), .S0 (nx4531)) ;
    xnor2 ix4634 (.Y (nx4633), .A0 (nx4635), .A1 (nx4637)) ;
    nand02 ix4636 (.Y (nx4635), .A0 (nx290), .A1 (nx5516)) ;
    xnor2 ix4638 (.Y (nx4637), .A0 (nx4639), .A1 (nx4641)) ;
    mux21 ix4640 (.Y (nx4639), .A0 (nx4537), .A1 (nx4543), .S0 (nx4539)) ;
    xnor2 ix4642 (.Y (nx4641), .A0 (nx4643), .A1 (nx4645)) ;
    nand02 ix4644 (.Y (nx4643), .A0 (nx266), .A1 (nx5512)) ;
    xnor2 ix4646 (.Y (nx4645), .A0 (nx4647), .A1 (nx4649)) ;
    mux21 ix4648 (.Y (nx4647), .A0 (nx4545), .A1 (nx4551), .S0 (nx4547)) ;
    xnor2 ix4650 (.Y (nx4649), .A0 (nx4651), .A1 (nx4653)) ;
    nand02 ix4652 (.Y (nx4651), .A0 (nx242), .A1 (nx5508)) ;
    xnor2 ix4654 (.Y (nx4653), .A0 (nx4655), .A1 (nx4657)) ;
    mux21 ix4656 (.Y (nx4655), .A0 (nx4553), .A1 (nx4559), .S0 (nx4555)) ;
    xnor2 ix4658 (.Y (nx4657), .A0 (nx4659), .A1 (nx4661)) ;
    nand02 ix4660 (.Y (nx4659), .A0 (nx218), .A1 (nx5504)) ;
    xnor2 ix4662 (.Y (nx4661), .A0 (nx4663), .A1 (nx4665)) ;
    mux21 ix4664 (.Y (nx4663), .A0 (nx4561), .A1 (nx4567), .S0 (nx4563)) ;
    xnor2 ix4666 (.Y (nx4665), .A0 (nx4667), .A1 (nx4669)) ;
    nand02 ix4668 (.Y (nx4667), .A0 (nx5500), .A1 (nx194)) ;
    xnor2 ix4670 (.Y (nx4669), .A0 (nx4671), .A1 (nx4673)) ;
    mux21 ix4672 (.Y (nx4671), .A0 (nx4569), .A1 (nx4575), .S0 (nx4571)) ;
    xnor2 ix4674 (.Y (nx4673), .A0 (nx4675), .A1 (nx4677)) ;
    nand02 ix4676 (.Y (nx4675), .A0 (nx5496), .A1 (nx170)) ;
    xnor2 ix4678 (.Y (nx4677), .A0 (nx4679), .A1 (nx4681)) ;
    mux21 ix4680 (.Y (nx4679), .A0 (nx4577), .A1 (nx4583), .S0 (nx4579)) ;
    xnor2 ix4682 (.Y (nx4681), .A0 (nx4683), .A1 (nx4685)) ;
    nand02 ix4684 (.Y (nx4683), .A0 (nx5492), .A1 (nx146)) ;
    xnor2 ix4686 (.Y (nx4685), .A0 (nx4687), .A1 (nx4689)) ;
    mux21 ix4688 (.Y (nx4687), .A0 (nx4585), .A1 (nx4591), .S0 (nx4587)) ;
    xnor2 ix4690 (.Y (nx4689), .A0 (nx4691), .A1 (nx4693)) ;
    nand02 ix4692 (.Y (nx4691), .A0 (nx5488), .A1 (nx122)) ;
    xnor2 ix4694 (.Y (nx4693), .A0 (nx4695), .A1 (nx4697)) ;
    mux21 ix4696 (.Y (nx4695), .A0 (nx4593), .A1 (nx4599), .S0 (nx4595)) ;
    xnor2 ix4698 (.Y (nx4697), .A0 (nx4699), .A1 (nx4701)) ;
    mux21 ix4702 (.Y (nx4701), .A0 (nx4601), .A1 (nx4607), .S0 (nx4603)) ;
    mux21 ix4704 (.Y (nx4703), .A0 (nx4519), .A1 (nx4609), .S0 (nx1903)) ;
    nor02 ix4475 (.Y (mac_output[22]), .A0 (RST), .A1 (nx4707)) ;
    nand02 ix4708 (.Y (nx4707), .A0 (nx2523), .A1 (nx4124)) ;
    xnor2 ix4125 (.Y (nx4124), .A0 (nx1901), .A1 (nx4789)) ;
    xnor2 ix4133 (.Y (nx1901), .A0 (mac_unit_tempP_22), .A1 (nx4714)) ;
    dffr mac_unit_MR_reg_Q_22 (.Q (mac_unit_tempP_22), .QB (\$dummy [53]), .D (
         nx4124), .CLK (CLK), .R (RST)) ;
    xnor2 ix4715 (.Y (nx4714), .A0 (nx4716), .A1 (nx4719)) ;
    mux21 ix4717 (.Y (nx4716), .A0 (nx4623), .A1 (nx4629), .S0 (nx4625)) ;
    xnor2 ix4720 (.Y (nx4719), .A0 (nx4721), .A1 (nx4723)) ;
    nand02 ix4722 (.Y (nx4721), .A0 (nx290), .A1 (nx5520)) ;
    xnor2 ix4724 (.Y (nx4723), .A0 (nx4725), .A1 (nx4727)) ;
    mux21 ix4726 (.Y (nx4725), .A0 (nx4631), .A1 (nx4637), .S0 (nx4633)) ;
    xnor2 ix4728 (.Y (nx4727), .A0 (nx4729), .A1 (nx4731)) ;
    nand02 ix4730 (.Y (nx4729), .A0 (nx266), .A1 (nx5516)) ;
    xnor2 ix4732 (.Y (nx4731), .A0 (nx4733), .A1 (nx4735)) ;
    mux21 ix4734 (.Y (nx4733), .A0 (nx4639), .A1 (nx4645), .S0 (nx4641)) ;
    xnor2 ix4736 (.Y (nx4735), .A0 (nx4737), .A1 (nx4739)) ;
    nand02 ix4738 (.Y (nx4737), .A0 (nx242), .A1 (nx5512)) ;
    xnor2 ix4740 (.Y (nx4739), .A0 (nx4741), .A1 (nx4743)) ;
    mux21 ix4742 (.Y (nx4741), .A0 (nx4647), .A1 (nx4653), .S0 (nx4649)) ;
    xnor2 ix4744 (.Y (nx4743), .A0 (nx4745), .A1 (nx4747)) ;
    nand02 ix4746 (.Y (nx4745), .A0 (nx218), .A1 (nx5508)) ;
    xnor2 ix4748 (.Y (nx4747), .A0 (nx4749), .A1 (nx4751)) ;
    mux21 ix4750 (.Y (nx4749), .A0 (nx4655), .A1 (nx4661), .S0 (nx4657)) ;
    xnor2 ix4752 (.Y (nx4751), .A0 (nx4753), .A1 (nx4755)) ;
    nand02 ix4754 (.Y (nx4753), .A0 (nx5504), .A1 (nx194)) ;
    xnor2 ix4756 (.Y (nx4755), .A0 (nx4757), .A1 (nx4759)) ;
    mux21 ix4758 (.Y (nx4757), .A0 (nx4663), .A1 (nx4669), .S0 (nx4665)) ;
    xnor2 ix4760 (.Y (nx4759), .A0 (nx4761), .A1 (nx4763)) ;
    nand02 ix4762 (.Y (nx4761), .A0 (nx5500), .A1 (nx170)) ;
    xnor2 ix4764 (.Y (nx4763), .A0 (nx4765), .A1 (nx4767)) ;
    mux21 ix4766 (.Y (nx4765), .A0 (nx4671), .A1 (nx4677), .S0 (nx4673)) ;
    xnor2 ix4768 (.Y (nx4767), .A0 (nx4769), .A1 (nx4771)) ;
    nand02 ix4770 (.Y (nx4769), .A0 (nx5496), .A1 (nx146)) ;
    xnor2 ix4772 (.Y (nx4771), .A0 (nx4773), .A1 (nx4775)) ;
    mux21 ix4774 (.Y (nx4773), .A0 (nx4679), .A1 (nx4685), .S0 (nx4681)) ;
    xnor2 ix4776 (.Y (nx4775), .A0 (nx4777), .A1 (nx4779)) ;
    nand02 ix4778 (.Y (nx4777), .A0 (nx5492), .A1 (nx122)) ;
    xnor2 ix4780 (.Y (nx4779), .A0 (nx4781), .A1 (nx4783)) ;
    mux21 ix4782 (.Y (nx4781), .A0 (nx4687), .A1 (nx4693), .S0 (nx4689)) ;
    xnor2 ix4784 (.Y (nx4783), .A0 (nx4785), .A1 (nx4787)) ;
    mux21 ix4788 (.Y (nx4787), .A0 (nx4695), .A1 (nx4701), .S0 (nx4697)) ;
    mux21 ix4790 (.Y (nx4789), .A0 (nx4620), .A1 (nx4703), .S0 (nx1902)) ;
    nor02 ix4483 (.Y (mac_output[23]), .A0 (RST), .A1 (nx4793)) ;
    nand02 ix4794 (.Y (nx4793), .A0 (nx2523), .A1 (nx4142)) ;
    xnor2 ix4143 (.Y (nx4142), .A0 (nx1899), .A1 (nx4865)) ;
    xnor2 ix4151 (.Y (nx1899), .A0 (mac_unit_tempP_23), .A1 (nx4799)) ;
    dffr mac_unit_MR_reg_Q_23 (.Q (mac_unit_tempP_23), .QB (\$dummy [54]), .D (
         nx4142), .CLK (CLK), .R (RST)) ;
    xnor2 ix4800 (.Y (nx4799), .A0 (nx4801), .A1 (nx4803)) ;
    mux21 ix4802 (.Y (nx4801), .A0 (nx4716), .A1 (nx4723), .S0 (nx4719)) ;
    xnor2 ix4804 (.Y (nx4803), .A0 (nx4805), .A1 (nx4807)) ;
    nand02 ix4806 (.Y (nx4805), .A0 (nx266), .A1 (nx5520)) ;
    xnor2 ix4808 (.Y (nx4807), .A0 (nx4809), .A1 (nx4811)) ;
    mux21 ix4810 (.Y (nx4809), .A0 (nx4725), .A1 (nx4731), .S0 (nx4727)) ;
    xnor2 ix4812 (.Y (nx4811), .A0 (nx4813), .A1 (nx4815)) ;
    nand02 ix4814 (.Y (nx4813), .A0 (nx242), .A1 (nx5516)) ;
    xnor2 ix4816 (.Y (nx4815), .A0 (nx4817), .A1 (nx4819)) ;
    mux21 ix4818 (.Y (nx4817), .A0 (nx4733), .A1 (nx4739), .S0 (nx4735)) ;
    xnor2 ix4820 (.Y (nx4819), .A0 (nx4821), .A1 (nx4823)) ;
    nand02 ix4822 (.Y (nx4821), .A0 (nx218), .A1 (nx5512)) ;
    xnor2 ix4824 (.Y (nx4823), .A0 (nx4825), .A1 (nx4827)) ;
    mux21 ix4826 (.Y (nx4825), .A0 (nx4741), .A1 (nx4747), .S0 (nx4743)) ;
    xnor2 ix4828 (.Y (nx4827), .A0 (nx4829), .A1 (nx4831)) ;
    nand02 ix4830 (.Y (nx4829), .A0 (nx194), .A1 (nx5508)) ;
    xnor2 ix4832 (.Y (nx4831), .A0 (nx4833), .A1 (nx4835)) ;
    mux21 ix4834 (.Y (nx4833), .A0 (nx4749), .A1 (nx4755), .S0 (nx4751)) ;
    xnor2 ix4836 (.Y (nx4835), .A0 (nx4837), .A1 (nx4839)) ;
    nand02 ix4838 (.Y (nx4837), .A0 (nx5504), .A1 (nx170)) ;
    xnor2 ix4840 (.Y (nx4839), .A0 (nx4841), .A1 (nx4843)) ;
    mux21 ix4842 (.Y (nx4841), .A0 (nx4757), .A1 (nx4763), .S0 (nx4759)) ;
    xnor2 ix4844 (.Y (nx4843), .A0 (nx4845), .A1 (nx4847)) ;
    nand02 ix4846 (.Y (nx4845), .A0 (nx5500), .A1 (nx146)) ;
    xnor2 ix4848 (.Y (nx4847), .A0 (nx4849), .A1 (nx4851)) ;
    mux21 ix4850 (.Y (nx4849), .A0 (nx4765), .A1 (nx4771), .S0 (nx4767)) ;
    xnor2 ix4852 (.Y (nx4851), .A0 (nx4853), .A1 (nx4855)) ;
    nand02 ix4854 (.Y (nx4853), .A0 (nx5496), .A1 (nx122)) ;
    xnor2 ix4856 (.Y (nx4855), .A0 (nx4857), .A1 (nx4859)) ;
    mux21 ix4858 (.Y (nx4857), .A0 (nx4773), .A1 (nx4779), .S0 (nx4775)) ;
    xnor2 ix4860 (.Y (nx4859), .A0 (nx4861), .A1 (nx4863)) ;
    mux21 ix4864 (.Y (nx4863), .A0 (nx4781), .A1 (nx4787), .S0 (nx4783)) ;
    mux21 ix4866 (.Y (nx4865), .A0 (nx4714), .A1 (nx4789), .S0 (nx1901)) ;
    nor02 ix4491 (.Y (mac_output[24]), .A0 (RST), .A1 (nx4868)) ;
    nand02 ix4869 (.Y (nx4868), .A0 (nx2523), .A1 (nx4160)) ;
    xnor2 ix4161 (.Y (nx4160), .A0 (nx1897), .A1 (nx4933)) ;
    xnor2 ix4169 (.Y (nx1897), .A0 (mac_unit_tempP_24), .A1 (nx4875)) ;
    dffr mac_unit_MR_reg_Q_24 (.Q (mac_unit_tempP_24), .QB (\$dummy [55]), .D (
         nx4160), .CLK (CLK), .R (RST)) ;
    xnor2 ix4876 (.Y (nx4875), .A0 (nx4877), .A1 (nx4879)) ;
    mux21 ix4878 (.Y (nx4877), .A0 (nx4801), .A1 (nx4807), .S0 (nx4803)) ;
    xnor2 ix4880 (.Y (nx4879), .A0 (nx4881), .A1 (nx4883)) ;
    nand02 ix4882 (.Y (nx4881), .A0 (nx242), .A1 (nx5520)) ;
    xnor2 ix4884 (.Y (nx4883), .A0 (nx4885), .A1 (nx4887)) ;
    mux21 ix4886 (.Y (nx4885), .A0 (nx4809), .A1 (nx4815), .S0 (nx4811)) ;
    xnor2 ix4888 (.Y (nx4887), .A0 (nx4889), .A1 (nx4891)) ;
    nand02 ix4890 (.Y (nx4889), .A0 (nx218), .A1 (nx5516)) ;
    xnor2 ix4892 (.Y (nx4891), .A0 (nx4893), .A1 (nx4895)) ;
    mux21 ix4894 (.Y (nx4893), .A0 (nx4817), .A1 (nx4823), .S0 (nx4819)) ;
    xnor2 ix4896 (.Y (nx4895), .A0 (nx4897), .A1 (nx4899)) ;
    nand02 ix4898 (.Y (nx4897), .A0 (nx194), .A1 (nx5512)) ;
    xnor2 ix4900 (.Y (nx4899), .A0 (nx4901), .A1 (nx4903)) ;
    mux21 ix4902 (.Y (nx4901), .A0 (nx4825), .A1 (nx4831), .S0 (nx4827)) ;
    xnor2 ix4904 (.Y (nx4903), .A0 (nx4905), .A1 (nx4907)) ;
    nand02 ix4906 (.Y (nx4905), .A0 (nx5508), .A1 (nx170)) ;
    xnor2 ix4908 (.Y (nx4907), .A0 (nx4909), .A1 (nx4911)) ;
    mux21 ix4910 (.Y (nx4909), .A0 (nx4833), .A1 (nx4839), .S0 (nx4835)) ;
    xnor2 ix4912 (.Y (nx4911), .A0 (nx4913), .A1 (nx4915)) ;
    nand02 ix4914 (.Y (nx4913), .A0 (nx5504), .A1 (nx146)) ;
    xnor2 ix4916 (.Y (nx4915), .A0 (nx4917), .A1 (nx4919)) ;
    mux21 ix4918 (.Y (nx4917), .A0 (nx4841), .A1 (nx4847), .S0 (nx4843)) ;
    xnor2 ix4920 (.Y (nx4919), .A0 (nx4921), .A1 (nx4923)) ;
    nand02 ix4922 (.Y (nx4921), .A0 (nx5500), .A1 (nx122)) ;
    xnor2 ix4924 (.Y (nx4923), .A0 (nx4925), .A1 (nx4927)) ;
    mux21 ix4926 (.Y (nx4925), .A0 (nx4849), .A1 (nx4855), .S0 (nx4851)) ;
    xnor2 ix4928 (.Y (nx4927), .A0 (nx4929), .A1 (nx4931)) ;
    mux21 ix4932 (.Y (nx4931), .A0 (nx4857), .A1 (nx4863), .S0 (nx4859)) ;
    mux21 ix4934 (.Y (nx4933), .A0 (nx4799), .A1 (nx4865), .S0 (nx1899)) ;
    nor02 ix4499 (.Y (mac_output[25]), .A0 (RST), .A1 (nx4937)) ;
    nand02 ix4938 (.Y (nx4937), .A0 (nx2523), .A1 (nx4178)) ;
    xnor2 ix4179 (.Y (nx4178), .A0 (nx1895), .A1 (nx4993)) ;
    xnor2 ix4187 (.Y (nx1895), .A0 (mac_unit_tempP_25), .A1 (nx4943)) ;
    dffr mac_unit_MR_reg_Q_25 (.Q (mac_unit_tempP_25), .QB (\$dummy [56]), .D (
         nx4178), .CLK (CLK), .R (RST)) ;
    xnor2 ix4944 (.Y (nx4943), .A0 (nx4945), .A1 (nx4947)) ;
    mux21 ix4946 (.Y (nx4945), .A0 (nx4877), .A1 (nx4883), .S0 (nx4879)) ;
    xnor2 ix4948 (.Y (nx4947), .A0 (nx4949), .A1 (nx4951)) ;
    nand02 ix4950 (.Y (nx4949), .A0 (nx218), .A1 (nx5520)) ;
    xnor2 ix4952 (.Y (nx4951), .A0 (nx4953), .A1 (nx4955)) ;
    mux21 ix4954 (.Y (nx4953), .A0 (nx4885), .A1 (nx4891), .S0 (nx4887)) ;
    xnor2 ix4956 (.Y (nx4955), .A0 (nx4957), .A1 (nx4959)) ;
    nand02 ix4958 (.Y (nx4957), .A0 (nx194), .A1 (nx5516)) ;
    xnor2 ix4960 (.Y (nx4959), .A0 (nx4961), .A1 (nx4963)) ;
    mux21 ix4962 (.Y (nx4961), .A0 (nx4893), .A1 (nx4899), .S0 (nx4895)) ;
    xnor2 ix4964 (.Y (nx4963), .A0 (nx4965), .A1 (nx4967)) ;
    nand02 ix4966 (.Y (nx4965), .A0 (nx170), .A1 (nx5512)) ;
    xnor2 ix4968 (.Y (nx4967), .A0 (nx4969), .A1 (nx4971)) ;
    mux21 ix4970 (.Y (nx4969), .A0 (nx4901), .A1 (nx4907), .S0 (nx4903)) ;
    xnor2 ix4972 (.Y (nx4971), .A0 (nx4973), .A1 (nx4975)) ;
    nand02 ix4974 (.Y (nx4973), .A0 (nx5508), .A1 (nx146)) ;
    xnor2 ix4976 (.Y (nx4975), .A0 (nx4977), .A1 (nx4979)) ;
    mux21 ix4978 (.Y (nx4977), .A0 (nx4909), .A1 (nx4915), .S0 (nx4911)) ;
    xnor2 ix4980 (.Y (nx4979), .A0 (nx4981), .A1 (nx4983)) ;
    nand02 ix4982 (.Y (nx4981), .A0 (nx5504), .A1 (nx122)) ;
    xnor2 ix4984 (.Y (nx4983), .A0 (nx4985), .A1 (nx4987)) ;
    mux21 ix4986 (.Y (nx4985), .A0 (nx4917), .A1 (nx4923), .S0 (nx4919)) ;
    xnor2 ix4988 (.Y (nx4987), .A0 (nx4989), .A1 (nx4991)) ;
    mux21 ix4992 (.Y (nx4991), .A0 (nx4925), .A1 (nx4931), .S0 (nx4927)) ;
    mux21 ix4994 (.Y (nx4993), .A0 (nx4875), .A1 (nx4933), .S0 (nx1897)) ;
    nor02 ix4507 (.Y (mac_output[26]), .A0 (RST), .A1 (nx4996)) ;
    nand02 ix4997 (.Y (nx4996), .A0 (nx2523), .A1 (nx4196)) ;
    xnor2 ix4197 (.Y (nx4196), .A0 (nx1893), .A1 (nx5044)) ;
    xnor2 ix4205 (.Y (nx1893), .A0 (mac_unit_tempP_26), .A1 (nx5002)) ;
    dffr mac_unit_MR_reg_Q_26 (.Q (mac_unit_tempP_26), .QB (\$dummy [57]), .D (
         nx4196), .CLK (CLK), .R (RST)) ;
    xnor2 ix5003 (.Y (nx5002), .A0 (nx5004), .A1 (nx5006)) ;
    mux21 ix5005 (.Y (nx5004), .A0 (nx4945), .A1 (nx4951), .S0 (nx4947)) ;
    xnor2 ix5007 (.Y (nx5006), .A0 (nx5008), .A1 (nx5010)) ;
    nand02 ix5009 (.Y (nx5008), .A0 (nx194), .A1 (nx5520)) ;
    xnor2 ix5011 (.Y (nx5010), .A0 (nx5012), .A1 (nx5014)) ;
    mux21 ix5013 (.Y (nx5012), .A0 (nx4953), .A1 (nx4959), .S0 (nx4955)) ;
    xnor2 ix5015 (.Y (nx5014), .A0 (nx5016), .A1 (nx5018)) ;
    nand02 ix5017 (.Y (nx5016), .A0 (nx170), .A1 (nx5516)) ;
    xnor2 ix5019 (.Y (nx5018), .A0 (nx5020), .A1 (nx5022)) ;
    mux21 ix5021 (.Y (nx5020), .A0 (nx4961), .A1 (nx4967), .S0 (nx4963)) ;
    xnor2 ix5023 (.Y (nx5022), .A0 (nx5024), .A1 (nx5026)) ;
    nand02 ix5025 (.Y (nx5024), .A0 (nx5512), .A1 (nx146)) ;
    xnor2 ix5027 (.Y (nx5026), .A0 (nx5028), .A1 (nx5030)) ;
    mux21 ix5029 (.Y (nx5028), .A0 (nx4969), .A1 (nx4975), .S0 (nx4971)) ;
    xnor2 ix5031 (.Y (nx5030), .A0 (nx5032), .A1 (nx5034)) ;
    nand02 ix5033 (.Y (nx5032), .A0 (nx5508), .A1 (nx122)) ;
    xnor2 ix5035 (.Y (nx5034), .A0 (nx5036), .A1 (nx5038)) ;
    mux21 ix5037 (.Y (nx5036), .A0 (nx4977), .A1 (nx4983), .S0 (nx4979)) ;
    xnor2 ix5039 (.Y (nx5038), .A0 (nx5040), .A1 (nx5042)) ;
    mux21 ix5043 (.Y (nx5042), .A0 (nx4985), .A1 (nx4991), .S0 (nx4987)) ;
    mux21 ix5045 (.Y (nx5044), .A0 (nx4943), .A1 (nx4993), .S0 (nx1895)) ;
    nor02 ix4515 (.Y (mac_output[27]), .A0 (RST), .A1 (nx5047)) ;
    nand02 ix5048 (.Y (nx5047), .A0 (nx2523), .A1 (nx4214)) ;
    xnor2 ix4215 (.Y (nx4214), .A0 (nx1892), .A1 (nx5087)) ;
    xnor2 ix4223 (.Y (nx1892), .A0 (mac_unit_tempP_27), .A1 (nx5053)) ;
    dffr mac_unit_MR_reg_Q_27 (.Q (mac_unit_tempP_27), .QB (\$dummy [58]), .D (
         nx4214), .CLK (CLK), .R (RST)) ;
    xnor2 ix5054 (.Y (nx5053), .A0 (nx5055), .A1 (nx5057)) ;
    mux21 ix5056 (.Y (nx5055), .A0 (nx5004), .A1 (nx5010), .S0 (nx5006)) ;
    xnor2 ix5058 (.Y (nx5057), .A0 (nx5059), .A1 (nx5061)) ;
    nand02 ix5060 (.Y (nx5059), .A0 (nx170), .A1 (nx5520)) ;
    xnor2 ix5062 (.Y (nx5061), .A0 (nx5063), .A1 (nx5065)) ;
    mux21 ix5064 (.Y (nx5063), .A0 (nx5012), .A1 (nx5018), .S0 (nx5014)) ;
    xnor2 ix5066 (.Y (nx5065), .A0 (nx5067), .A1 (nx5069)) ;
    nand02 ix5068 (.Y (nx5067), .A0 (nx146), .A1 (nx5516)) ;
    xnor2 ix5070 (.Y (nx5069), .A0 (nx5071), .A1 (nx5073)) ;
    mux21 ix5072 (.Y (nx5071), .A0 (nx5020), .A1 (nx5026), .S0 (nx5022)) ;
    xnor2 ix5074 (.Y (nx5073), .A0 (nx5075), .A1 (nx5077)) ;
    nand02 ix5076 (.Y (nx5075), .A0 (nx5512), .A1 (nx122)) ;
    xnor2 ix5078 (.Y (nx5077), .A0 (nx5079), .A1 (nx5081)) ;
    mux21 ix5080 (.Y (nx5079), .A0 (nx5028), .A1 (nx5034), .S0 (nx5030)) ;
    xnor2 ix5082 (.Y (nx5081), .A0 (nx5083), .A1 (nx5085)) ;
    mux21 ix5086 (.Y (nx5085), .A0 (nx5036), .A1 (nx5042), .S0 (nx5038)) ;
    mux21 ix5088 (.Y (nx5087), .A0 (nx5002), .A1 (nx5044), .S0 (nx1893)) ;
    nor02 ix4523 (.Y (mac_output[28]), .A0 (RST), .A1 (nx5090)) ;
    nand02 ix5091 (.Y (nx5090), .A0 (nx2523), .A1 (nx4232)) ;
    xnor2 ix4233 (.Y (nx4232), .A0 (nx1891), .A1 (nx5122)) ;
    xnor2 ix4241 (.Y (nx1891), .A0 (mac_unit_tempP_28), .A1 (nx5096)) ;
    dffr mac_unit_MR_reg_Q_28 (.Q (mac_unit_tempP_28), .QB (\$dummy [59]), .D (
         nx4232), .CLK (CLK), .R (RST)) ;
    xnor2 ix5097 (.Y (nx5096), .A0 (nx5098), .A1 (nx5100)) ;
    mux21 ix5099 (.Y (nx5098), .A0 (nx5055), .A1 (nx5061), .S0 (nx5057)) ;
    xnor2 ix5101 (.Y (nx5100), .A0 (nx5102), .A1 (nx5104)) ;
    nand02 ix5103 (.Y (nx5102), .A0 (nx146), .A1 (nx5520)) ;
    xnor2 ix5105 (.Y (nx5104), .A0 (nx5106), .A1 (nx5108)) ;
    mux21 ix5107 (.Y (nx5106), .A0 (nx5063), .A1 (nx5069), .S0 (nx5065)) ;
    xnor2 ix5109 (.Y (nx5108), .A0 (nx5110), .A1 (nx5112)) ;
    nand02 ix5111 (.Y (nx5110), .A0 (nx5516), .A1 (nx122)) ;
    xnor2 ix5113 (.Y (nx5112), .A0 (nx5114), .A1 (nx5116)) ;
    mux21 ix5115 (.Y (nx5114), .A0 (nx5071), .A1 (nx5077), .S0 (nx5073)) ;
    xnor2 ix5117 (.Y (nx5116), .A0 (nx5118), .A1 (nx5120)) ;
    mux21 ix5121 (.Y (nx5120), .A0 (nx5079), .A1 (nx5085), .S0 (nx5081)) ;
    mux21 ix5123 (.Y (nx5122), .A0 (nx5053), .A1 (nx5087), .S0 (nx1892)) ;
    nor02 ix4531 (.Y (mac_output[29]), .A0 (RST), .A1 (nx5125)) ;
    nand02 ix5126 (.Y (nx5125), .A0 (nx2523), .A1 (nx4250)) ;
    xnor2 ix4251 (.Y (nx4250), .A0 (nx1889), .A1 (nx5149)) ;
    xnor2 ix4259 (.Y (nx1889), .A0 (mac_unit_tempP_29), .A1 (nx5131)) ;
    dffr mac_unit_MR_reg_Q_29 (.Q (mac_unit_tempP_29), .QB (\$dummy [60]), .D (
         nx4250), .CLK (CLK), .R (RST)) ;
    xnor2 ix5132 (.Y (nx5131), .A0 (nx5133), .A1 (nx5135)) ;
    mux21 ix5134 (.Y (nx5133), .A0 (nx5098), .A1 (nx5104), .S0 (nx5100)) ;
    xnor2 ix5136 (.Y (nx5135), .A0 (nx5137), .A1 (nx5139)) ;
    nand02 ix5138 (.Y (nx5137), .A0 (nx122), .A1 (nx5520)) ;
    xnor2 ix5140 (.Y (nx5139), .A0 (nx5141), .A1 (nx5143)) ;
    mux21 ix5142 (.Y (nx5141), .A0 (nx5106), .A1 (nx5112), .S0 (nx5108)) ;
    xnor2 ix5144 (.Y (nx5143), .A0 (nx5145), .A1 (nx5147)) ;
    mux21 ix5148 (.Y (nx5147), .A0 (nx5114), .A1 (nx5120), .S0 (nx5116)) ;
    mux21 ix5150 (.Y (nx5149), .A0 (nx5096), .A1 (nx5122), .S0 (nx1891)) ;
    nor02 ix4539 (.Y (mac_output[30]), .A0 (RST), .A1 (nx5152)) ;
    nand02 ix5153 (.Y (nx5152), .A0 (nx2523), .A1 (nx4268)) ;
    xnor2 ix4269 (.Y (nx4268), .A0 (nx1887), .A1 (nx5168)) ;
    xnor2 ix4277 (.Y (nx1887), .A0 (mac_unit_tempP_30), .A1 (nx5158)) ;
    dffr mac_unit_MR_reg_Q_30 (.Q (mac_unit_tempP_30), .QB (\$dummy [61]), .D (
         nx4268), .CLK (CLK), .R (RST)) ;
    xnor2 ix5159 (.Y (nx5158), .A0 (nx5160), .A1 (nx5162)) ;
    mux21 ix5161 (.Y (nx5160), .A0 (nx5133), .A1 (nx5139), .S0 (nx5135)) ;
    xnor2 ix5163 (.Y (nx5162), .A0 (nx5164), .A1 (nx5166)) ;
    mux21 ix5167 (.Y (nx5166), .A0 (nx5141), .A1 (nx5147), .S0 (nx5143)) ;
    mux21 ix5169 (.Y (nx5168), .A0 (nx5131), .A1 (nx5149), .S0 (nx1889)) ;
    nor02ii ix4291 (.Y (mac_output[31]), .A0 (RST), .A1 (nx1885)) ;
    xnor2 ix4287 (.Y (nx1885), .A0 (nx3636), .A1 (nx5177)) ;
    xnor2 ix3637 (.Y (nx3636), .A0 (mac_unit_tempP_31), .A1 (nx5175)) ;
    dffr mac_unit_MR_reg_Q_31 (.Q (mac_unit_tempP_31), .QB (\$dummy [62]), .D (
         nx1885), .CLK (CLK), .R (RST)) ;
    mux21 ix5176 (.Y (nx5175), .A0 (nx5160), .A1 (nx5166), .S0 (nx5162)) ;
    mux21 ix5178 (.Y (nx5177), .A0 (nx5158), .A1 (nx5168), .S0 (nx1887)) ;
    dff test_output_reg_signature_0 (.Q (sig_0), .QB (\$dummy [63]), .D (
        test_output_misr_signal_31), .CLK (CLK)) ;
    oai32 ix2416 (.Y (nx2415), .A0 (nx5183), .A1 (RST), .A2 (nx5526), .B0 (
          nx5345), .B1 (nx5542)) ;
    xnor2 ix5184 (.Y (nx5183), .A0 (nx4294), .A1 (test_output_misr_signal_30)) ;
    nor02 ix4295 (.Y (nx4294), .A0 (RST), .A1 (nx2429)) ;
    dffr test_output_reg_misr_signal_30 (.Q (test_output_misr_signal_30), .QB (
         \$dummy [64]), .D (nx2405), .CLK (CLK), .R (RST)) ;
    oai32 ix2396 (.Y (nx2395), .A0 (nx5191), .A1 (RST), .A2 (nx5526), .B0 (
          nx5342), .B1 (nx5542)) ;
    oai32 ix2386 (.Y (nx2385), .A0 (nx5195), .A1 (RST), .A2 (nx5526), .B0 (
          nx5340), .B1 (nx5542)) ;
    oai32 ix2376 (.Y (nx2375), .A0 (nx5199), .A1 (RST), .A2 (nx5526), .B0 (
          nx5338), .B1 (nx5542)) ;
    oai32 ix2366 (.Y (nx2365), .A0 (nx5203), .A1 (RST), .A2 (nx5526), .B0 (
          nx5336), .B1 (nx5542)) ;
    oai32 ix2356 (.Y (nx2355), .A0 (nx5207), .A1 (RST), .A2 (nx5526), .B0 (
          nx5334), .B1 (nx5446)) ;
    oai32 ix2346 (.Y (nx2345), .A0 (nx5211), .A1 (RST), .A2 (nx5526), .B0 (
          nx5332), .B1 (nx5446)) ;
    oai32 ix2336 (.Y (nx2335), .A0 (nx5215), .A1 (RST), .A2 (nx5524), .B0 (
          nx5330), .B1 (nx5446)) ;
    oai32 ix2326 (.Y (nx2325), .A0 (nx5219), .A1 (RST), .A2 (nx5524), .B0 (
          nx5328), .B1 (nx5446)) ;
    oai32 ix2316 (.Y (nx2315), .A0 (nx5223), .A1 (RST), .A2 (nx5524), .B0 (
          nx5326), .B1 (nx5446)) ;
    oai32 ix2306 (.Y (nx2305), .A0 (nx5227), .A1 (RST), .A2 (nx5524), .B0 (
          nx5324), .B1 (nx5446)) ;
    oai32 ix2296 (.Y (nx2295), .A0 (nx5231), .A1 (RST), .A2 (nx5524), .B0 (
          nx5322), .B1 (nx5446)) ;
    oai32 ix2286 (.Y (nx2285), .A0 (nx5235), .A1 (RST), .A2 (nx5524), .B0 (
          nx5320), .B1 (nx5446)) ;
    oai32 ix2276 (.Y (nx2275), .A0 (nx5239), .A1 (RST), .A2 (nx5524), .B0 (
          nx5318), .B1 (nx5446)) ;
    oai32 ix2266 (.Y (nx2265), .A0 (nx5243), .A1 (RST), .A2 (nx5524), .B0 (
          nx5316), .B1 (nx5446)) ;
    oai32 ix2256 (.Y (nx2255), .A0 (nx5247), .A1 (RST), .A2 (nx5524), .B0 (
          nx5314), .B1 (nx5446)) ;
    xnor2 ix5248 (.Y (nx5247), .A0 (nx4422), .A1 (test_output_misr_signal_14)) ;
    dffr test_output_reg_misr_signal_14 (.Q (test_output_misr_signal_14), .QB (
         \$dummy [65]), .D (nx2245), .CLK (CLK), .R (RST)) ;
    oai32 ix2236 (.Y (nx2235), .A0 (nx5254), .A1 (RST), .A2 (nx5524), .B0 (
          nx5311), .B1 (nx5446)) ;
    xnor2 ix5255 (.Y (nx5254), .A0 (nx4438), .A1 (test_output_misr_signal_12)) ;
    dffr test_output_reg_misr_signal_12 (.Q (test_output_misr_signal_12), .QB (
         \$dummy [66]), .D (nx2225), .CLK (CLK), .R (RST)) ;
    xnor2 ix4617 (.Y (nx4616), .A0 (nx4391), .A1 (test_output_misr_signal_11)) ;
    dffr test_output_reg_misr_signal_11 (.Q (test_output_misr_signal_11), .QB (
         \$dummy [67]), .D (nx2215), .CLK (CLK), .R (RST)) ;
    xnor2 ix4611 (.Y (nx4610), .A0 (nx4511), .A1 (test_output_misr_signal_10)) ;
    dffr test_output_reg_misr_signal_10 (.Q (test_output_misr_signal_10), .QB (
         \$dummy [68]), .D (nx2205), .CLK (CLK), .R (RST)) ;
    xnor2 ix4605 (.Y (nx4604), .A0 (nx4613), .A1 (test_output_misr_signal_9)) ;
    dffr test_output_reg_misr_signal_9 (.Q (test_output_misr_signal_9), .QB (
         \$dummy [69]), .D (nx2195), .CLK (CLK), .R (RST)) ;
    xnor2 ix4599 (.Y (nx4598), .A0 (nx4707), .A1 (test_output_misr_signal_8)) ;
    dffr test_output_reg_misr_signal_8 (.Q (test_output_misr_signal_8), .QB (
         \$dummy [70]), .D (nx2185), .CLK (CLK), .R (RST)) ;
    xnor2 ix4593 (.Y (nx4592), .A0 (nx4793), .A1 (test_output_misr_signal_7)) ;
    dffr test_output_reg_misr_signal_7 (.Q (test_output_misr_signal_7), .QB (
         \$dummy [71]), .D (nx2175), .CLK (CLK), .R (RST)) ;
    xnor2 ix4587 (.Y (nx4586), .A0 (nx4868), .A1 (test_output_misr_signal_6)) ;
    dffr test_output_reg_misr_signal_6 (.Q (test_output_misr_signal_6), .QB (
         \$dummy [72]), .D (nx2165), .CLK (CLK), .R (RST)) ;
    xnor2 ix4581 (.Y (nx4580), .A0 (nx4937), .A1 (test_output_misr_signal_5)) ;
    dffr test_output_reg_misr_signal_5 (.Q (test_output_misr_signal_5), .QB (
         \$dummy [73]), .D (nx2155), .CLK (CLK), .R (RST)) ;
    xnor2 ix4575 (.Y (nx4574), .A0 (nx4996), .A1 (test_output_misr_signal_4)) ;
    dffr test_output_reg_misr_signal_4 (.Q (test_output_misr_signal_4), .QB (
         \$dummy [74]), .D (nx2145), .CLK (CLK), .R (RST)) ;
    xnor2 ix4569 (.Y (nx4568), .A0 (nx5047), .A1 (test_output_misr_signal_3)) ;
    dffr test_output_reg_misr_signal_3 (.Q (test_output_misr_signal_3), .QB (
         \$dummy [75]), .D (nx2135), .CLK (CLK), .R (RST)) ;
    xnor2 ix4563 (.Y (nx4562), .A0 (nx5090), .A1 (test_output_misr_signal_2)) ;
    dffr test_output_reg_misr_signal_2 (.Q (test_output_misr_signal_2), .QB (
         \$dummy [76]), .D (nx2125), .CLK (CLK), .R (RST)) ;
    xnor2 ix4557 (.Y (nx4556), .A0 (nx5125), .A1 (test_output_misr_signal_1)) ;
    dffr test_output_reg_misr_signal_1 (.Q (test_output_misr_signal_1), .QB (
         \$dummy [77]), .D (nx2115), .CLK (CLK), .R (RST)) ;
    xnor2 ix4551 (.Y (nx4550), .A0 (nx5152), .A1 (test_output_misr_signal_0)) ;
    dffr test_output_reg_misr_signal_0 (.Q (test_output_misr_signal_0), .QB (
         \$dummy [78]), .D (nx2105), .CLK (CLK), .R (RST)) ;
    xnor2 ix4545 (.Y (nx4544), .A0 (nx4868), .A1 (nx4542)) ;
    dffr test_output_reg_misr_signal_13 (.Q (test_output_misr_signal_13), .QB (
         nx5311), .D (nx2235), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_15 (.Q (test_output_misr_signal_15), .QB (
         nx5314), .D (nx2255), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_16 (.Q (test_output_misr_signal_16), .QB (
         nx5316), .D (nx2265), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_17 (.Q (test_output_misr_signal_17), .QB (
         nx5318), .D (nx2275), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_18 (.Q (test_output_misr_signal_18), .QB (
         nx5320), .D (nx2285), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_19 (.Q (test_output_misr_signal_19), .QB (
         nx5322), .D (nx2295), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_20 (.Q (test_output_misr_signal_20), .QB (
         nx5324), .D (nx2305), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_21 (.Q (test_output_misr_signal_21), .QB (
         nx5326), .D (nx2315), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_22 (.Q (test_output_misr_signal_22), .QB (
         nx5328), .D (nx2325), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_23 (.Q (test_output_misr_signal_23), .QB (
         nx5330), .D (nx2335), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_24 (.Q (test_output_misr_signal_24), .QB (
         nx5332), .D (nx2345), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_25 (.Q (test_output_misr_signal_25), .QB (
         nx5334), .D (nx2355), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_26 (.Q (test_output_misr_signal_26), .QB (
         nx5336), .D (nx2365), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_27 (.Q (test_output_misr_signal_27), .QB (
         nx5338), .D (nx2375), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_28 (.Q (test_output_misr_signal_28), .QB (
         nx5340), .D (nx2385), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_29 (.Q (test_output_misr_signal_29), .QB (
         nx5342), .D (nx2395), .CLK (CLK), .R (RST)) ;
    dffr test_output_reg_misr_signal_31 (.Q (test_output_misr_signal_31), .QB (
         nx5345), .D (nx2415), .CLK (CLK), .R (RST)) ;
    dff test_output_reg_signature_1 (.Q (sig_1), .QB (\$dummy [79]), .D (
        test_output_misr_signal_30), .CLK (CLK)) ;
    dff test_output_reg_signature_2 (.Q (sig_2), .QB (\$dummy [80]), .D (
        test_output_misr_signal_29), .CLK (CLK)) ;
    dff test_output_reg_signature_3 (.Q (sig_3), .QB (\$dummy [81]), .D (
        test_output_misr_signal_28), .CLK (CLK)) ;
    dff test_output_reg_signature_4 (.Q (sig_4), .QB (\$dummy [82]), .D (
        test_output_misr_signal_27), .CLK (CLK)) ;
    dff test_output_reg_signature_5 (.Q (sig_5), .QB (\$dummy [83]), .D (
        test_output_misr_signal_26), .CLK (CLK)) ;
    dff test_output_reg_signature_6 (.Q (sig_6), .QB (\$dummy [84]), .D (
        test_output_misr_signal_25), .CLK (CLK)) ;
    dff test_output_reg_signature_7 (.Q (sig_7), .QB (\$dummy [85]), .D (
        test_output_misr_signal_24), .CLK (CLK)) ;
    dff test_output_reg_signature_8 (.Q (sig_8), .QB (\$dummy [86]), .D (
        test_output_misr_signal_23), .CLK (CLK)) ;
    dff test_output_reg_signature_9 (.Q (sig_9), .QB (\$dummy [87]), .D (
        test_output_misr_signal_22), .CLK (CLK)) ;
    dff test_output_reg_signature_10 (.Q (sig_10), .QB (\$dummy [88]), .D (
        test_output_misr_signal_21), .CLK (CLK)) ;
    dff test_output_reg_signature_11 (.Q (sig_11), .QB (\$dummy [89]), .D (
        test_output_misr_signal_20), .CLK (CLK)) ;
    dff test_output_reg_signature_12 (.Q (sig_12), .QB (\$dummy [90]), .D (
        test_output_misr_signal_19), .CLK (CLK)) ;
    dff test_output_reg_signature_13 (.Q (sig_13), .QB (\$dummy [91]), .D (
        test_output_misr_signal_18), .CLK (CLK)) ;
    dff test_output_reg_signature_14 (.Q (sig_14), .QB (\$dummy [92]), .D (
        test_output_misr_signal_17), .CLK (CLK)) ;
    dff test_output_reg_signature_15 (.Q (sig_15), .QB (\$dummy [93]), .D (
        test_output_misr_signal_16), .CLK (CLK)) ;
    dff test_output_reg_signature_16 (.Q (sig_16), .QB (\$dummy [94]), .D (
        test_output_misr_signal_15), .CLK (CLK)) ;
    dff test_output_reg_signature_17 (.Q (sig_17), .QB (\$dummy [95]), .D (
        test_output_misr_signal_14), .CLK (CLK)) ;
    dff test_output_reg_signature_18 (.Q (sig_18), .QB (\$dummy [96]), .D (
        test_output_misr_signal_13), .CLK (CLK)) ;
    dff test_output_reg_signature_19 (.Q (sig_19), .QB (\$dummy [97]), .D (
        test_output_misr_signal_12), .CLK (CLK)) ;
    dff test_output_reg_signature_20 (.Q (sig_20), .QB (\$dummy [98]), .D (
        test_output_misr_signal_11), .CLK (CLK)) ;
    dff test_output_reg_signature_21 (.Q (sig_21), .QB (\$dummy [99]), .D (
        test_output_misr_signal_10), .CLK (CLK)) ;
    dff test_output_reg_signature_22 (.Q (sig_22), .QB (\$dummy [100]), .D (
        test_output_misr_signal_9), .CLK (CLK)) ;
    dff test_output_reg_signature_23 (.Q (sig_23), .QB (\$dummy [101]), .D (
        test_output_misr_signal_8), .CLK (CLK)) ;
    dff test_output_reg_signature_24 (.Q (sig_24), .QB (\$dummy [102]), .D (
        test_output_misr_signal_7), .CLK (CLK)) ;
    dff test_output_reg_signature_25 (.Q (sig_25), .QB (\$dummy [103]), .D (
        test_output_misr_signal_6), .CLK (CLK)) ;
    dff test_output_reg_signature_26 (.Q (sig_26), .QB (\$dummy [104]), .D (
        test_output_misr_signal_5), .CLK (CLK)) ;
    dff test_output_reg_signature_27 (.Q (sig_27), .QB (\$dummy [105]), .D (
        test_output_misr_signal_4), .CLK (CLK)) ;
    dff test_output_reg_signature_28 (.Q (sig_28), .QB (\$dummy [106]), .D (
        test_output_misr_signal_3), .CLK (CLK)) ;
    dff test_output_reg_signature_29 (.Q (sig_29), .QB (\$dummy [107]), .D (
        test_output_misr_signal_2), .CLK (CLK)) ;
    dff test_output_reg_signature_30 (.Q (sig_30), .QB (\$dummy [108]), .D (
        test_output_misr_signal_1), .CLK (CLK)) ;
    dff test_output_reg_signature_31 (.Q (sig_31), .QB (\$dummy [109]), .D (
        test_output_misr_signal_0), .CLK (CLK)) ;
    inv01 ix4053 (.Y (nx4052), .A (nx4251)) ;
    inv01 ix4051 (.Y (nx4050), .A (nx4257)) ;
    inv01 ix4017 (.Y (nx4016), .A (nx3963)) ;
    inv01 ix4015 (.Y (nx4014), .A (nx3971)) ;
    inv01 ix3993 (.Y (nx3992), .A (nx3815)) ;
    inv01 ix3991 (.Y (nx3990), .A (nx3823)) ;
    inv01 ix3969 (.Y (nx3968), .A (nx3681)) ;
    inv01 ix3967 (.Y (nx3966), .A (nx3687)) ;
    inv01 ix3945 (.Y (nx3944), .A (nx3549)) ;
    inv01 ix3943 (.Y (nx3942), .A (nx3557)) ;
    inv01 ix3921 (.Y (nx3920), .A (nx3425)) ;
    inv01 ix3919 (.Y (nx3918), .A (nx3433)) ;
    inv01 ix3897 (.Y (nx3896), .A (nx3311)) ;
    inv01 ix3895 (.Y (nx3894), .A (nx3319)) ;
    inv01 ix3873 (.Y (nx3872), .A (nx3203)) ;
    inv01 ix3871 (.Y (nx3870), .A (nx3211)) ;
    inv01 ix3849 (.Y (nx3848), .A (nx3103)) ;
    inv01 ix3847 (.Y (nx3846), .A (nx3111)) ;
    inv01 ix3825 (.Y (nx3824), .A (nx3011)) ;
    inv01 ix3823 (.Y (nx3822), .A (nx3019)) ;
    inv01 ix3801 (.Y (nx3800), .A (nx2921)) ;
    inv01 ix3799 (.Y (nx3798), .A (nx2929)) ;
    inv01 ix3777 (.Y (nx3776), .A (nx2839)) ;
    inv01 ix3775 (.Y (nx3774), .A (nx2847)) ;
    inv01 ix3753 (.Y (nx3752), .A (nx2765)) ;
    inv01 ix3751 (.Y (nx3750), .A (nx2773)) ;
    inv01 ix3729 (.Y (nx3728), .A (nx2699)) ;
    inv01 ix3727 (.Y (nx3726), .A (nx2707)) ;
    inv01 ix3705 (.Y (nx3704), .A (nx2643)) ;
    inv01 ix3703 (.Y (nx3702), .A (nx2651)) ;
    inv01 ix3681 (.Y (nx3680), .A (nx2601)) ;
    inv01 ix3679 (.Y (nx3678), .A (nx2609)) ;
    inv01 ix3639 (.Y (nx3638), .A (nx2429)) ;
    inv01 ix3695 (.Y (nx1933), .A (nx2603)) ;
    inv01 ix3719 (.Y (nx1932), .A (nx2645)) ;
    inv01 ix3743 (.Y (nx1931), .A (nx2701)) ;
    inv01 ix3767 (.Y (nx1929), .A (nx2767)) ;
    inv01 ix3791 (.Y (nx1927), .A (nx2841)) ;
    inv01 ix3815 (.Y (nx1925), .A (nx2923)) ;
    inv01 ix3839 (.Y (nx1923), .A (nx3013)) ;
    inv01 ix3863 (.Y (nx1922), .A (nx3105)) ;
    inv01 ix3887 (.Y (nx1921), .A (nx3205)) ;
    inv01 ix3911 (.Y (nx1919), .A (nx3313)) ;
    inv01 ix3935 (.Y (nx1917), .A (nx3427)) ;
    inv01 ix3959 (.Y (nx1915), .A (nx3551)) ;
    inv01 ix3983 (.Y (nx1913), .A (nx3683)) ;
    inv01 ix4007 (.Y (nx1912), .A (nx3817)) ;
    inv01 ix4025 (.Y (nx1911), .A (nx3965)) ;
    inv01 ix4061 (.Y (nx1907), .A (nx4253)) ;
    inv01 ix4110 (.Y (nx4109), .A (nx3574)) ;
    inv01 ix4404 (.Y (nx4403), .A (nx3540)) ;
    inv01 ix3956 (.Y (nx3955), .A (nx3420)) ;
    inv01 ix4414 (.Y (nx4413), .A (nx3364)) ;
    inv01 ix3808 (.Y (nx3807), .A (nx3198)) ;
    inv01 ix3996 (.Y (nx3995), .A (nx3134)) ;
    inv01 ix4128 (.Y (nx4127), .A (nx3096)) ;
    inv01 ix4280 (.Y (nx4279), .A (nx3086)) ;
    inv01 ix3674 (.Y (nx3673), .A (nx2976)) ;
    inv01 ix3856 (.Y (nx3855), .A (nx2912)) ;
    inv01 ix4138 (.Y (nx4137), .A (nx2864)) ;
    inv01 ix4290 (.Y (nx4289), .A (nx2854)) ;
    inv01 ix3542 (.Y (nx3541), .A (nx2754)) ;
    inv01 ix3718 (.Y (nx3717), .A (nx2690)) ;
    inv01 ix4148 (.Y (nx4147), .A (nx2632)) ;
    inv01 ix4300 (.Y (nx4299), .A (nx2622)) ;
    inv01 ix3418 (.Y (nx3417), .A (nx2532)) ;
    inv01 ix3590 (.Y (nx3589), .A (nx2468)) ;
    inv01 ix4158 (.Y (nx4157), .A (nx2400)) ;
    inv01 ix4310 (.Y (nx4309), .A (nx2390)) ;
    inv01 ix3304 (.Y (nx3303), .A (nx2310)) ;
    inv01 ix3466 (.Y (nx3465), .A (nx2246)) ;
    inv01 ix4168 (.Y (nx4167), .A (nx2168)) ;
    inv01 ix4320 (.Y (nx4319), .A (nx2158)) ;
    inv01 ix3196 (.Y (nx3195), .A (nx2088)) ;
    inv01 ix3352 (.Y (nx3351), .A (nx2024)) ;
    inv01 ix4178 (.Y (nx4177), .A (nx1936)) ;
    inv01 ix4330 (.Y (nx4329), .A (nx1926)) ;
    inv01 ix3096 (.Y (nx3095), .A (nx1866)) ;
    inv01 ix3244 (.Y (nx3243), .A (nx1802)) ;
    inv01 ix4188 (.Y (nx4187), .A (nx1704)) ;
    inv01 ix4340 (.Y (nx4339), .A (nx1694)) ;
    inv01 ix3004 (.Y (nx3003), .A (nx1644)) ;
    inv01 ix3144 (.Y (nx3143), .A (nx1580)) ;
    inv01 ix4198 (.Y (nx4197), .A (nx1472)) ;
    inv01 ix4350 (.Y (nx4349), .A (nx1462)) ;
    inv01 ix2914 (.Y (nx2913), .A (nx1422)) ;
    inv01 ix3052 (.Y (nx3051), .A (nx1358)) ;
    inv01 ix4206 (.Y (nx4205), .A (nx1240)) ;
    inv01 ix4360 (.Y (nx4359), .A (nx1230)) ;
    inv01 ix2832 (.Y (nx2831), .A (nx1200)) ;
    inv01 ix2966 (.Y (nx2965), .A (nx1136)) ;
    inv01 ix4216 (.Y (nx4215), .A (nx1008)) ;
    inv01 ix4370 (.Y (nx4369), .A (nx998)) ;
    inv01 ix2758 (.Y (nx2757), .A (nx978)) ;
    inv01 ix2884 (.Y (nx2883), .A (nx914)) ;
    inv01 ix4224 (.Y (nx4223), .A (nx776)) ;
    inv01 ix4380 (.Y (nx4379), .A (nx766)) ;
    inv01 ix2692 (.Y (nx2691), .A (nx756)) ;
    inv01 ix2810 (.Y (nx2809), .A (nx692)) ;
    inv01 ix4234 (.Y (nx4233), .A (nx544)) ;
    inv01 ix2636 (.Y (nx2635), .A (nx528)) ;
    inv01 ix4388 (.Y (nx4387), .A (nx520)) ;
    inv01 ix2744 (.Y (nx2743), .A (nx464)) ;
    inv01 ix2580 (.Y (nx2579), .A (nx456)) ;
    inv01 ix2592 (.Y (nx2591), .A (nx434)) ;
    inv01 ix2584 (.Y (nx2583), .A (nx114)) ;
    inv01 ix4092 (.Y (nx4091), .A (nx98)) ;
    inv01 ix2588 (.Y (nx2587), .A (nx90)) ;
    inv01 ix5445 (.Y (nx5446), .A (nx5534)) ;
    inv01 ix5447 (.Y (nx5448), .A (nx2587)) ;
    inv01 ix5449 (.Y (nx5450), .A (nx2587)) ;
    inv01 ix5455 (.Y (nx5456), .A (nx2583)) ;
    inv01 ix5463 (.Y (nx5464), .A (nx5548)) ;
    inv01 ix5467 (.Y (nx5468), .A (nx2635)) ;
    inv01 ix5471 (.Y (nx5472), .A (nx2691)) ;
    inv01 ix5475 (.Y (nx5476), .A (nx2757)) ;
    inv01 ix5479 (.Y (nx5480), .A (nx2831)) ;
    inv01 ix5483 (.Y (nx5484), .A (nx2913)) ;
    inv01 ix5487 (.Y (nx5488), .A (nx3003)) ;
    inv01 ix5491 (.Y (nx5492), .A (nx3095)) ;
    inv01 ix5495 (.Y (nx5496), .A (nx3195)) ;
    inv01 ix5499 (.Y (nx5500), .A (nx3303)) ;
    inv01 ix5503 (.Y (nx5504), .A (nx3417)) ;
    inv01 ix5507 (.Y (nx5508), .A (nx3541)) ;
    inv01 ix5511 (.Y (nx5512), .A (nx3673)) ;
    inv01 ix5515 (.Y (nx5516), .A (nx3807)) ;
    inv01 ix5519 (.Y (nx5520), .A (nx3955)) ;
    inv01 ix5523 (.Y (nx5524), .A (test_mode)) ;
    inv01 ix5525 (.Y (nx5526), .A (test_mode)) ;
    inv02 ix5533 (.Y (nx5534), .A (nx10)) ;
    inv01 ix5535 (.Y (nx5536), .A (nx456)) ;
    or02 ix2440 (.Y (nx2439), .A0 (nx2587), .A1 (nx5548)) ;
    mux21 ix2096 (.Y (nx2095), .A0 (test_input_lfsr_signal_15), .A1 (
          test_input_lfsr_signal_14), .S0 (nx5542)) ;
    mux21 ix2086 (.Y (nx2085), .A0 (test_input_lfsr_signal_14), .A1 (
          test_input_lfsr_signal_13), .S0 (nx5542)) ;
    mux21 ix2076 (.Y (nx2075), .A0 (test_input_lfsr_signal_13), .A1 (
          test_input_lfsr_signal_12), .S0 (nx5542)) ;
    mux21 ix2066 (.Y (nx2065), .A0 (test_input_lfsr_signal_12), .A1 (
          test_input_lfsr_signal_11), .S0 (nx5542)) ;
    mux21 ix2056 (.Y (nx2055), .A0 (test_input_lfsr_signal_11), .A1 (
          test_input_lfsr_signal_10), .S0 (nx5542)) ;
    mux21 ix2046 (.Y (nx2045), .A0 (test_input_lfsr_signal_10), .A1 (
          test_input_lfsr_signal_9), .S0 (nx5542)) ;
    mux21 ix2036 (.Y (nx2035), .A0 (test_input_lfsr_signal_9), .A1 (
          test_input_lfsr_signal_8), .S0 (nx5542)) ;
    mux21 ix2026 (.Y (nx2025), .A0 (test_input_lfsr_signal_8), .A1 (
          test_input_lfsr_signal_7), .S0 (nx5542)) ;
    mux21 ix2016 (.Y (nx2015), .A0 (test_input_lfsr_signal_7), .A1 (
          test_input_lfsr_signal_6), .S0 (nx5542)) ;
    mux21 ix2006 (.Y (nx2005), .A0 (test_input_lfsr_signal_6), .A1 (
          test_input_lfsr_signal_5), .S0 (nx5542)) ;
    mux21 ix1996 (.Y (nx1995), .A0 (test_input_lfsr_signal_5), .A1 (
          test_input_lfsr_signal_4), .S0 (nx5544)) ;
    mux21 ix1986 (.Y (nx1985), .A0 (test_input_lfsr_signal_4), .A1 (
          test_input_lfsr_signal_3), .S0 (nx5544)) ;
    mux21 ix1976 (.Y (nx1975), .A0 (test_input_lfsr_signal_3), .A1 (
          test_input_lfsr_signal_2), .S0 (nx5544)) ;
    mux21 ix1966 (.Y (nx1965), .A0 (test_input_lfsr_signal_2), .A1 (
          test_input_lfsr_signal_1), .S0 (nx5544)) ;
    mux21 ix1956 (.Y (nx1955), .A0 (test_input_lfsr_signal_1), .A1 (
          test_input_lfsr_signal_0), .S0 (nx5544)) ;
    nor02ii ix2522 (.Y (nx10), .A0 (RST), .A1 (test_mode)) ;
    or04 ix2568 (.Y (nx2567), .A0 (nx2587), .A1 (nx5548), .A2 (nx2583), .A3 (
         nx2591)) ;
    ao22 ix3665 (.Y (nx3664), .A0 (nx456), .A1 (nx114), .B0 (nx90), .B1 (nx434)
         ) ;
    or02 ix2614 (.Y (nx2613), .A0 (nx5548), .A1 (nx2635)) ;
    or02 ix2626 (.Y (nx2625), .A0 (nx2583), .A1 (nx2591)) ;
    or02 ix2662 (.Y (nx2661), .A0 (nx5548), .A1 (nx2691)) ;
    or02 ix2674 (.Y (nx2673), .A0 (nx2591), .A1 (nx2635)) ;
    or02 ix2718 (.Y (nx2717), .A0 (nx5548), .A1 (nx2757)) ;
    or02 ix2730 (.Y (nx2729), .A0 (nx2591), .A1 (nx2691)) ;
    or02 ix2784 (.Y (nx2783), .A0 (nx5548), .A1 (nx2831)) ;
    or02 ix2796 (.Y (nx2795), .A0 (nx2591), .A1 (nx2757)) ;
    or02 ix2858 (.Y (nx2857), .A0 (nx5548), .A1 (nx2913)) ;
    or02 ix2870 (.Y (nx2869), .A0 (nx2591), .A1 (nx2831)) ;
    or02 ix2940 (.Y (nx2939), .A0 (nx5548), .A1 (nx3003)) ;
    or02 ix2952 (.Y (nx2951), .A0 (nx2591), .A1 (nx2913)) ;
    or02 ix3030 (.Y (nx3029), .A0 (nx5548), .A1 (nx3095)) ;
    or02 ix3038 (.Y (nx3037), .A0 (nx2591), .A1 (nx3003)) ;
    or02 ix3122 (.Y (nx3121), .A0 (nx5548), .A1 (nx3195)) ;
    or02 ix3130 (.Y (nx3129), .A0 (nx2591), .A1 (nx3095)) ;
    or02 ix3222 (.Y (nx3221), .A0 (nx5548), .A1 (nx3303)) ;
    or02 ix3230 (.Y (nx3229), .A0 (nx2591), .A1 (nx3195)) ;
    or02 ix3330 (.Y (nx3329), .A0 (nx5548), .A1 (nx3417)) ;
    or02 ix3338 (.Y (nx3337), .A0 (nx2591), .A1 (nx3303)) ;
    or02 ix3444 (.Y (nx3443), .A0 (nx5548), .A1 (nx3541)) ;
    or02 ix3452 (.Y (nx3451), .A0 (nx2591), .A1 (nx3417)) ;
    or02 ix3568 (.Y (nx3567), .A0 (nx5548), .A1 (nx3673)) ;
    or02 ix3576 (.Y (nx3575), .A0 (nx2591), .A1 (nx3541)) ;
    or02 ix3698 (.Y (nx3697), .A0 (nx2579), .A1 (nx3807)) ;
    or02 ix3706 (.Y (nx3705), .A0 (nx2591), .A1 (nx3673)) ;
    or02 ix3834 (.Y (nx3833), .A0 (nx2579), .A1 (nx3955)) ;
    or02 ix3842 (.Y (nx3841), .A0 (nx2591), .A1 (nx3807)) ;
    or02 ix3950 (.Y (nx3949), .A0 (nx2587), .A1 (nx5550)) ;
    or02 ix3982 (.Y (nx3981), .A0 (nx2591), .A1 (nx3955)) ;
    or02 ix4086 (.Y (nx4085), .A0 (nx2583), .A1 (nx5550)) ;
    or02 ix4238 (.Y (nx4237), .A0 (nx2635), .A1 (nx5550)) ;
    or02 ix4384 (.Y (nx4383), .A0 (nx2691), .A1 (nx5550)) ;
    or02 ix4498 (.Y (nx4497), .A0 (nx2757), .A1 (nx5550)) ;
    or02 ix4606 (.Y (nx4605), .A0 (nx2831), .A1 (nx5550)) ;
    or02 ix4700 (.Y (nx4699), .A0 (nx2913), .A1 (nx5550)) ;
    or02 ix4786 (.Y (nx4785), .A0 (nx3003), .A1 (nx5550)) ;
    or02 ix4862 (.Y (nx4861), .A0 (nx3095), .A1 (nx5550)) ;
    or02 ix4930 (.Y (nx4929), .A0 (nx3195), .A1 (nx5550)) ;
    or02 ix4990 (.Y (nx4989), .A0 (nx3303), .A1 (nx5550)) ;
    or02 ix5041 (.Y (nx5040), .A0 (nx3417), .A1 (nx5550)) ;
    or02 ix5084 (.Y (nx5083), .A0 (nx3541), .A1 (nx5550)) ;
    or02 ix5119 (.Y (nx5118), .A0 (nx3673), .A1 (nx5550)) ;
    or02 ix5146 (.Y (nx5145), .A0 (nx3807), .A1 (nx4091)) ;
    or02 ix5165 (.Y (nx5164), .A0 (nx3955), .A1 (nx4091)) ;
    and02 ix4743 (.Y (signature[0]), .A0 (test_mode), .A1 (sig_0)) ;
    mux21 ix2406 (.Y (nx2405), .A0 (test_output_misr_signal_30), .A1 (nx4724), .S0 (
          nx5544)) ;
    xor2 ix4725 (.Y (nx4724), .A0 (nx2555), .A1 (nx5342)) ;
    xor2 ix5192 (.Y (nx5191), .A0 (nx4310), .A1 (nx5340)) ;
    xor2 ix5196 (.Y (nx5195), .A0 (nx4318), .A1 (nx5338)) ;
    xor2 ix5200 (.Y (nx5199), .A0 (nx4326), .A1 (nx5336)) ;
    xor2 ix5204 (.Y (nx5203), .A0 (nx4334), .A1 (nx5334)) ;
    xor2 ix5208 (.Y (nx5207), .A0 (nx4342), .A1 (nx5332)) ;
    xor2 ix5212 (.Y (nx5211), .A0 (nx4350), .A1 (nx5330)) ;
    xor2 ix5216 (.Y (nx5215), .A0 (nx4358), .A1 (nx5328)) ;
    xor2 ix5220 (.Y (nx5219), .A0 (nx4366), .A1 (nx5326)) ;
    xor2 ix5224 (.Y (nx5223), .A0 (nx4374), .A1 (nx5324)) ;
    xor2 ix5228 (.Y (nx5227), .A0 (nx4382), .A1 (nx5322)) ;
    xor2 ix5232 (.Y (nx5231), .A0 (nx4390), .A1 (nx5320)) ;
    xor2 ix5236 (.Y (nx5235), .A0 (nx4398), .A1 (nx5318)) ;
    xor2 ix5240 (.Y (nx5239), .A0 (nx4406), .A1 (nx5316)) ;
    xor2 ix5244 (.Y (nx5243), .A0 (nx4414), .A1 (nx5314)) ;
    mux21 ix2246 (.Y (nx2245), .A0 (test_output_misr_signal_14), .A1 (nx4628), .S0 (
          nx5544)) ;
    xor2 ix4629 (.Y (nx4628), .A0 (nx4095), .A1 (nx5311)) ;
    mux21 ix2226 (.Y (nx2225), .A0 (test_output_misr_signal_12), .A1 (nx4616), .S0 (
          nx5544)) ;
    mux21 ix2216 (.Y (nx2215), .A0 (test_output_misr_signal_11), .A1 (nx4610), .S0 (
          nx5544)) ;
    mux21 ix2206 (.Y (nx2205), .A0 (test_output_misr_signal_10), .A1 (nx4604), .S0 (
          nx5544)) ;
    mux21 ix2196 (.Y (nx2195), .A0 (test_output_misr_signal_9), .A1 (nx4598), .S0 (
          nx5544)) ;
    mux21 ix2186 (.Y (nx2185), .A0 (test_output_misr_signal_8), .A1 (nx4592), .S0 (
          nx5544)) ;
    mux21 ix2176 (.Y (nx2175), .A0 (test_output_misr_signal_7), .A1 (nx4586), .S0 (
          nx5544)) ;
    mux21 ix2166 (.Y (nx2165), .A0 (test_output_misr_signal_6), .A1 (nx4580), .S0 (
          nx5544)) ;
    mux21 ix2156 (.Y (nx2155), .A0 (test_output_misr_signal_5), .A1 (nx4574), .S0 (
          nx5544)) ;
    mux21 ix2146 (.Y (nx2145), .A0 (test_output_misr_signal_4), .A1 (nx4568), .S0 (
          nx5546)) ;
    mux21 ix2136 (.Y (nx2135), .A0 (test_output_misr_signal_3), .A1 (nx4562), .S0 (
          nx5546)) ;
    mux21 ix2126 (.Y (nx2125), .A0 (test_output_misr_signal_2), .A1 (nx4556), .S0 (
          nx5546)) ;
    mux21 ix2116 (.Y (nx2115), .A0 (test_output_misr_signal_1), .A1 (nx4550), .S0 (
          nx5546)) ;
    mux21 ix2106 (.Y (nx2105), .A0 (test_output_misr_signal_0), .A1 (nx4544), .S0 (
          nx5546)) ;
    xor2 ix4543 (.Y (nx4542), .A0 (nx5334), .A1 (nx5296)) ;
    xnor2 ix5297 (.Y (nx5296), .A0 (nx5345), .A1 (nx5342)) ;
    and02 ix4751 (.Y (signature[1]), .A0 (test_mode), .A1 (sig_1)) ;
    and02 ix4759 (.Y (signature[2]), .A0 (test_mode), .A1 (sig_2)) ;
    and02 ix4767 (.Y (signature[3]), .A0 (test_mode), .A1 (sig_3)) ;
    and02 ix4775 (.Y (signature[4]), .A0 (test_mode), .A1 (sig_4)) ;
    and02 ix4783 (.Y (signature[5]), .A0 (test_mode), .A1 (sig_5)) ;
    and02 ix4791 (.Y (signature[6]), .A0 (test_mode), .A1 (sig_6)) ;
    and02 ix4799 (.Y (signature[7]), .A0 (test_mode), .A1 (sig_7)) ;
    and02 ix4807 (.Y (signature[8]), .A0 (test_mode), .A1 (sig_8)) ;
    and02 ix4815 (.Y (signature[9]), .A0 (test_mode), .A1 (sig_9)) ;
    and02 ix4823 (.Y (signature[10]), .A0 (test_mode), .A1 (sig_10)) ;
    and02 ix4831 (.Y (signature[11]), .A0 (test_mode), .A1 (sig_11)) ;
    and02 ix4839 (.Y (signature[12]), .A0 (test_mode), .A1 (sig_12)) ;
    and02 ix4847 (.Y (signature[13]), .A0 (test_mode), .A1 (sig_13)) ;
    and02 ix4855 (.Y (signature[14]), .A0 (test_mode), .A1 (sig_14)) ;
    and02 ix4863 (.Y (signature[15]), .A0 (test_mode), .A1 (sig_15)) ;
    and02 ix4871 (.Y (signature[16]), .A0 (test_mode), .A1 (sig_16)) ;
    and02 ix4879 (.Y (signature[17]), .A0 (test_mode), .A1 (sig_17)) ;
    and02 ix4887 (.Y (signature[18]), .A0 (test_mode), .A1 (sig_18)) ;
    and02 ix4895 (.Y (signature[19]), .A0 (test_mode), .A1 (sig_19)) ;
    and02 ix4903 (.Y (signature[20]), .A0 (test_mode), .A1 (sig_20)) ;
    and02 ix4911 (.Y (signature[21]), .A0 (test_mode), .A1 (sig_21)) ;
    and02 ix4919 (.Y (signature[22]), .A0 (test_mode), .A1 (sig_22)) ;
    and02 ix4927 (.Y (signature[23]), .A0 (test_mode), .A1 (sig_23)) ;
    and02 ix4935 (.Y (signature[24]), .A0 (test_mode), .A1 (sig_24)) ;
    and02 ix4943 (.Y (signature[25]), .A0 (test_mode), .A1 (sig_25)) ;
    and02 ix4951 (.Y (signature[26]), .A0 (test_mode), .A1 (sig_26)) ;
    and02 ix4959 (.Y (signature[27]), .A0 (test_mode), .A1 (sig_27)) ;
    and02 ix4967 (.Y (signature[28]), .A0 (test_mode), .A1 (sig_28)) ;
    and02 ix4975 (.Y (signature[29]), .A0 (test_mode), .A1 (sig_29)) ;
    and02 ix4983 (.Y (signature[30]), .A0 (test_mode), .A1 (sig_30)) ;
    and02 ix4991 (.Y (signature[31]), .A0 (test_mode), .A1 (sig_31)) ;
    inv02 ix5541 (.Y (nx5542), .A (nx5534)) ;
    inv02 ix5543 (.Y (nx5544), .A (nx5534)) ;
    inv02 ix5545 (.Y (nx5546), .A (nx5534)) ;
    inv01 ix5547 (.Y (nx5548), .A (nx456)) ;
    inv01 ix5549 (.Y (nx5550), .A (nx98)) ;
endmodule

